`include "common.h"

module chip_z80(
  input eclk, ereset,
  output ab0,
  output ab1,
  output ab2,
  output ab3,
  output ab4,
  output ab5,
  output ab6,
  output ab7,
  output ab8,
  output ab9,
  output ab10,
  output ab11,
  output ab12,
  output ab13,
  output ab14,
  output ab15,
  input db0_i,
  output db0_o,
  output db0_t,
  input db1_i,
  output db1_o,
  output db1_t,
  input db2_i,
  output db2_o,
  output db2_t,
  input db3_i,
  output db3_o,
  output db3_t,
  input db4_i,
  output db4_o,
  output db4_t,
  input db5_i,
  output db5_o,
  output db5_t,
  input db6_i,
  output db6_o,
  output db6_t,
  input db7_i,
  output db7_o,
  output db7_t,
  input _reset,
  input _wait,
  input _int,
  input _nmi,
  input _busrq,
  output _m1,
  output _rd,
  output _wr,
  output _mreq,
  output _iorq,
  output _rfsh,
  output _halt,
  output _busak,
  input clk
);

  function v;   // convert an analog node value to 2-level
  input [`W-1:0] x;
  begin
    v = ~x[`W-1];
  end
  endfunction

  function [`W-1:0] a;   // convert a 2-level node value to analog
  input x;
  begin
    a = x ? `HI2 : `LO2;
  end
  endfunction

  wire signed [`W-1:0] n_779_port_3, n_779_port_4, n_779_port_5, n_779_port_8, n_779_v;
  wire signed [`W-1:0] n_791_port_0, n_791_port_1, n_791_port_3, n_791_port_4, n_791_v;
  wire signed [`W-1:0] n_1498_port_2, n_1498_port_3, n_1498_v;
  wire signed [`W-1:0] n_703_port_0, n_703_port_3, n_703_port_4, n_703_port_5, n_703_v;
  wire signed [`W-1:0] n_907_port_0, n_907_port_3, n_907_port_4, n_907_port_5, n_907_v;
  wire signed [`W-1:0] db0_port_0, db0_port_1, db0_port_3, db0_v;
  wire signed [`W-1:0] db7_port_0, db7_port_2, db7_port_3, db7_v;
  wire signed [`W-1:0] n_783_port_5, n_783_port_6, n_783_port_7, n_783_port_8, n_783_port_9, n_783_port_10, n_783_v;
  wire signed [`W-1:0] db1_port_0, db1_port_2, db1_port_3, db1_v;
  wire signed [`W-1:0] n_380_port_0, n_380_port_2, n_380_v;
  wire signed [`W-1:0] n_480_port_0, n_480_port_7, n_480_v;
  wire signed [`W-1:0] n_485_port_0, n_485_port_7, n_485_v;
  wire signed [`W-1:0] n_486_port_0, n_486_port_6, n_486_v;
  wire signed [`W-1:0] n_713_port_0, n_713_port_1, n_713_port_3, n_713_port_4, n_713_v;
  wire signed [`W-1:0] n_545_port_4, n_545_port_8, n_545_port_10, n_545_port_11, n_545_port_12, n_545_port_14, n_545_v;
  wire signed [`W-1:0] n_917_port_0, n_917_port_1, n_917_port_3, n_917_port_4, n_917_v;
  wire signed [`W-1:0] n_798_port_0, n_798_port_2, n_798_port_3, n_798_port_4, n_798_v;
  wire signed [`W-1:0] n_370_port_0, n_370_port_4, n_370_v;
  wire signed [`W-1:0] n_196_port_0, n_196_port_4, n_196_v;
  wire signed [`W-1:0] n_412_port_0, n_412_port_4, n_412_v;
  wire signed [`W-1:0] n_138_port_0, n_138_port_3, n_138_v;
  wire signed [`W-1:0] n_790_port_0, n_790_port_1, n_790_port_3, n_790_port_5, n_790_v;
  wire signed [`W-1:0] n_922_port_0, n_922_port_2, n_922_port_3, n_922_port_4, n_922_v;
  wire signed [`W-1:0] n_806_port_0, n_806_port_3, n_806_port_4, n_806_port_5, n_806_v;
  wire signed [`W-1:0] n_525_port_3, n_525_port_7, n_525_port_8, n_525_port_9, n_525_port_11, n_525_port_13, n_525_port_15, n_525_v;
  wire signed [`W-1:0] n_808_port_5, n_808_port_6, n_808_port_7, n_808_port_8, n_808_port_9, n_808_port_10, n_808_v;
  wire signed [`W-1:0] n_2338_port_0, n_2338_port_3, n_2338_port_5, n_2338_v;
  wire signed [`W-1:0] n_796_port_5, n_796_port_6, n_796_port_7, n_796_port_8, n_796_port_9, n_796_port_10, n_796_v;
  wire signed [`W-1:0] n_933_port_0, n_933_port_3, n_933_port_4, n_933_port_5, n_933_v;
  wire signed [`W-1:0] n_714_port_0, n_714_port_2, n_714_port_3, n_714_port_4, n_714_v;
  wire signed [`W-1:0] db6_port_0, db6_port_1, db6_port_3, db6_v;
  wire signed [`W-1:0] n_248_port_0, n_248_port_25, n_248_port_26, n_248_v;
  wire signed [`W-1:0] n_1332_port_1, n_1332_port_2, n_1332_v;
  wire signed [`W-1:0] n_73_port_4, n_73_port_6, n_73_v;
  wire signed [`W-1:0] n_528_port_0, n_528_port_1, n_528_port_3, n_528_port_6, n_528_port_7, n_528_v;
  wire signed [`W-1:0] n_810_port_0, n_810_port_3, n_810_port_4, n_810_port_5, n_810_v;
  wire signed [`W-1:0] n_936_port_0, n_936_port_3, n_936_port_4, n_936_port_5, n_936_v;
  wire signed [`W-1:0] n_731_port_0, n_731_port_3, n_731_port_4, n_731_port_5, n_731_v;
  wire signed [`W-1:0] n_616_port_0, n_616_port_1, n_616_v;
  wire signed [`W-1:0] n_803_port_5, n_803_port_6, n_803_port_7, n_803_port_8, n_803_port_9, n_803_port_10, n_803_v;
  wire signed [`W-1:0] n_944_port_0, n_944_port_2, n_944_port_3, n_944_port_4, n_944_v;
  wire signed [`W-1:0] n_716_port_0, n_716_port_3, n_716_port_4, n_716_port_7, n_716_port_8, n_716_v;
  wire signed [`W-1:0] n_947_port_0, n_947_port_2, n_947_port_3, n_947_port_4, n_947_v;
  wire signed [`W-1:0] n_953_port_0, n_953_port_1, n_953_port_3, n_953_port_4, n_953_v;
  wire signed [`W-1:0] n_841_port_0, n_841_port_1, n_841_port_3, n_841_port_4, n_841_v;
  wire signed [`W-1:0] db2_port_0, db2_port_1, db2_port_3, db2_v;
  wire signed [`W-1:0] n_845_port_0, n_845_port_2, n_845_port_3, n_845_port_4, n_845_v;
  wire signed [`W-1:0] n_958_port_0, n_958_port_2, n_958_port_3, n_958_port_4, n_958_v;
  wire signed [`W-1:0] n_755_port_5, n_755_port_6, n_755_port_7, n_755_port_8, n_755_port_9, n_755_v;
  wire signed [`W-1:0] n_846_port_0, n_846_port_2, n_846_port_3, n_846_port_4, n_846_v;
  wire signed [`W-1:0] n_739_port_0, n_739_port_3, n_739_port_4, n_739_port_5, n_739_v;
  wire signed [`W-1:0] n_850_port_0, n_850_port_2, n_850_port_3, n_850_port_4, n_850_v;
  wire signed [`W-1:0] n_969_port_0, n_969_port_3, n_969_port_4, n_969_port_5, n_969_v;
  wire signed [`W-1:0] n_863_port_0, n_863_port_3, n_863_port_4, n_863_port_5, n_863_v;
  wire signed [`W-1:0] db5_port_0, db5_port_1, db5_port_3, db5_v;
  wire signed [`W-1:0] n_526_port_0, n_526_port_3, n_526_port_6, n_526_port_7, n_526_port_8, n_526_v;
  wire signed [`W-1:0] db3_port_0, db3_port_2, db3_port_3, db3_v;
  wire signed [`W-1:0] n_749_port_0, n_749_port_1, n_749_port_3, n_749_port_4, n_749_v;
  wire signed [`W-1:0] n_974_port_0, n_974_port_3, n_974_port_4, n_974_port_5, n_974_v;
  wire signed [`W-1:0] n_836_port_5, n_836_port_6, n_836_port_7, n_836_port_8, n_836_port_9, n_836_port_10, n_836_v;
  wire signed [`W-1:0] n_2504_port_0, n_2504_port_3, n_2504_port_5, n_2504_v;
  wire signed [`W-1:0] n_966_port_0, n_966_port_2, n_966_port_3, n_966_port_4, n_966_v;
  wire signed [`W-1:0] n_982_port_0, n_982_port_1, n_982_port_3, n_982_port_4, n_982_v;
  wire signed [`W-1:0] n_681_port_5, n_681_port_6, n_681_port_7, n_681_port_8, n_681_port_9, n_681_v;
  wire signed [`W-1:0] n_871_port_0, n_871_port_3, n_871_port_4, n_871_port_5, n_871_v;
  wire signed [`W-1:0] n_752_port_0, n_752_port_2, n_752_port_3, n_752_port_4, n_752_v;
  wire signed [`W-1:0] n_984_port_0, n_984_port_2, n_984_port_3, n_984_port_4, n_984_v;
  wire signed [`W-1:0] n_562_v;
  wire signed [`W-1:0] n_993_port_0, n_993_port_2, n_993_port_3, n_993_port_4, n_993_v;
  wire signed [`W-1:0] n_839_port_5, n_839_port_6, n_839_port_7, n_839_port_8, n_839_port_9, n_839_v;
  wire signed [`W-1:0] n_2211_port_0, n_2211_port_3, n_2211_port_5, n_2211_v;
  wire signed [`W-1:0] n_884_port_0, n_884_port_1, n_884_port_3, n_884_port_4, n_884_v;
  wire signed [`W-1:0] n_998_port_0, n_998_port_3, n_998_port_4, n_998_port_5, n_998_v;
  wire signed [`W-1:0] n_770_port_2, n_770_port_4, n_770_port_5, n_770_port_6, n_770_v;
  wire signed [`W-1:0] n_774_port_0, n_774_port_3, n_774_port_4, n_774_port_5, n_774_v;
  wire signed [`W-1:0] n_885_port_0, n_885_port_2, n_885_port_3, n_885_port_4, n_885_v;
  wire signed [`W-1:0] n_816_port_0, n_816_port_4, n_816_port_6, n_816_v;
  wire signed [`W-1:0] n_1005_port_3, n_1005_port_4, n_1005_port_5, n_1005_port_6, n_1005_v;
  wire signed [`W-1:0] n_772_port_5, n_772_port_6, n_772_port_7, n_772_port_8, n_772_port_9, n_772_port_10, n_772_v;
  wire signed [`W-1:0] clk_port_403, clk_v;
  wire signed [`W-1:0] ex_bcdehl_port_5, ex_bcdehl_port_8, ex_bcdehl_v;
  wire signed [`W-1:0] n_897_port_0, n_897_port_2, n_897_port_3, n_897_port_4, n_897_v;
  wire signed [`W-1:0] n_901_port_0, n_901_port_2, n_901_port_3, n_901_port_5, n_901_v;
  wire signed [`W-1:0] n_899_port_0, n_899_port_2, n_899_port_3, n_899_port_4, n_899_v;
  wire signed [`W-1:0] n_697_port_0, n_697_port_1, n_697_port_3, n_697_port_4, n_697_port_5, n_697_v;
  wire signed [`W-1:0] n_777_port_0, n_777_port_3, n_777_port_4, n_777_port_5, n_777_v;
  wire signed [`W-1:0] n_124_port_5, n_124_port_9, n_124_v;
  wire signed [`W-1:0] n_45_v;
  wire signed [`W-1:0] db4_port_0, db4_port_1, db4_port_3, db4_v;
  wire signed [`W-1:0] n_175_port_3, n_175_port_6, n_175_v;
  wire signed [`W-1:0] n_1225_port_5, n_1225_port_7, n_1225_v;
  wire signed [`W-1:0] n_181_port_4, n_181_port_5, n_181_port_6, n_181_port_7, n_181_v;
  wire signed [`W-1:0] n_176_port_5, n_176_port_10, n_176_v;
  wire signed [`W-1:0] n_1232_port_3, n_1232_port_5, n_1232_v;
  wire signed [`W-1:0] n_190_port_0, n_190_port_3, n_190_v;
  wire signed [`W-1:0] n_1218_port_3, n_1218_port_6, n_1218_v;
  wire signed [`W-1:0] n_1228_port_5, n_1228_port_7, n_1228_v;
  wire signed [`W-1:0] n_1220_port_6, n_1220_port_10, n_1220_v;
  wire signed [`W-1:0] n_172_port_4, n_172_port_8, n_172_v;
  wire signed [`W-1:0] n_1168_port_4, n_1168_port_8, n_1168_v;
  wire signed [`W-1:0] n_1466_port_3, n_1466_port_4, n_1466_v;
  wire signed [`W-1:0] n_1161_port_4, n_1161_port_9, n_1161_v;
  wire signed [`W-1:0] n_1051_port_3, n_1051_port_6, n_1051_v;
  wire signed [`W-1:0] n_75_port_5, n_75_port_6, n_75_v;
  wire signed [`W-1:0] n_77_port_5, n_77_port_8, n_77_v;
  wire signed [`W-1:0] n_1060_port_3, n_1060_port_5, n_1060_v;
  wire signed [`W-1:0] n_185_port_5, n_185_port_7, n_185_v;
  wire signed [`W-1:0] n_61_port_3, n_61_port_5, n_61_v;
  wire signed [`W-1:0] n_1053_port_4, n_1053_port_6, n_1053_v;
  wire signed [`W-1:0] n_136_port_5, n_136_port_10, n_136_v;
  wire signed [`W-1:0] n_1221_port_5, n_1221_port_7, n_1221_v;
  wire signed [`W-1:0] _nmi_port_1, _nmi_v;
  wire signed [`W-1:0] n_56_port_5, n_56_port_11, n_56_v;
  wire signed [`W-1:0] n_1271_port_4, n_1271_port_6, n_1271_v;
  wire signed [`W-1:0] n_223_port_3, n_223_port_6, n_223_v;
  wire signed [`W-1:0] n_68_port_4, n_68_port_9, n_68_v;
  wire signed [`W-1:0] n_58_port_4, n_58_port_8, n_58_v;
  wire signed [`W-1:0] n_197_port_3, n_197_port_6, n_197_v;
  wire signed [`W-1:0] n_148_port_6, n_148_port_13, n_148_v;
  wire signed [`W-1:0] n_57_port_3, n_57_port_6, n_57_v;
  wire signed [`W-1:0] n_67_port_3, n_67_port_5, n_67_v;
  wire signed [`W-1:0] n_92_port_4, n_92_port_7, n_92_v;
  wire signed [`W-1:0] n_1092_port_3, n_1092_port_5, n_1092_v;
  wire signed [`W-1:0] n_1043_port_1, n_1043_port_3, n_1043_v;
  wire signed [`W-1:0] n_1080_port_4, n_1080_port_8, n_1080_v;
  wire signed [`W-1:0] n_1590_port_1, n_1590_port_2, n_1590_port_3, n_1590_v;
  wire signed [`W-1:0] n_1095_port_4, n_1095_port_8, n_1095_v;
  wire signed [`W-1:0] n_120_port_5, n_120_port_9, n_120_v;
  wire signed [`W-1:0] n_1079_port_3, n_1079_port_5, n_1079_v;
  wire signed [`W-1:0] n_128_port_6, n_128_port_10, n_128_v;
  wire signed [`W-1:0] n_1300_port_2, n_1300_port_3, n_1300_v;
  wire signed [`W-1:0] n_1302_port_0, n_1302_port_2, n_1302_v;
  wire signed [`W-1:0] n_1586_port_4, n_1586_port_6, n_1586_v;
  wire signed [`W-1:0] n_139_port_5, n_139_port_12, n_139_v;
  wire signed [`W-1:0] n_1126_port_5, n_1126_port_8, n_1126_v;
  wire signed [`W-1:0] n_70_port_4, n_70_port_7, n_70_v;
  wire signed [`W-1:0] _busrq_port_1, _busrq_v;
  wire signed [`W-1:0] _wait_port_1, _wait_v;
  wire signed [`W-1:0] n_241_port_5, n_241_port_7, n_241_v;
  wire signed [`W-1:0] n_216_port_5, n_216_port_8, n_216_v;
  wire signed [`W-1:0] n_1320_port_3, n_1320_port_5, n_1320_v;
  wire signed [`W-1:0] n_240_port_5, n_240_port_8, n_240_v;
  wire signed [`W-1:0] n_214_port_3, n_214_port_5, n_214_v;
  wire signed [`W-1:0] n_150_port_5, n_150_port_11, n_150_v;
  wire signed [`W-1:0] n_1313_port_3, n_1313_port_6, n_1313_v;
  wire signed [`W-1:0] n_1701_port_4, n_1701_port_8, n_1701_v;
  wire signed [`W-1:0] ex_dehl0_port_5, ex_dehl0_port_9, ex_dehl0_v;
  wire signed [`W-1:0] n_1702_port_4, n_1702_port_8, n_1702_v;
  wire signed [`W-1:0] ex_dehl1_port_5, ex_dehl1_port_9, ex_dehl1_v;
  wire signed [`W-1:0] n_1709_v;
  wire signed [`W-1:0] n_244_port_4, n_244_port_8, n_244_v;
  wire signed [`W-1:0] _int_port_1, _int_v;
  wire signed [`W-1:0] n_633_port_5, n_633_port_9, n_633_v;
  wire signed [`W-1:0] n_84_port_6, n_84_port_10, n_84_v;
  wire signed [`W-1:0] n_1129_port_3, n_1129_port_6, n_1129_v;
  wire signed [`W-1:0] ex_af_port_5, ex_af_port_10, ex_af_v;
  wire signed [`W-1:0] n_647_port_0, n_647_port_3, n_647_port_4, n_647_port_5, n_647_v;
  wire signed [`W-1:0] n_687_port_5, n_687_port_6, n_687_v;
  wire signed [`W-1:0] n_1783_port_4, n_1783_port_6, n_1783_v;
  wire signed [`W-1:0] n_1773_port_5, n_1773_port_9, n_1773_v;
  wire signed [`W-1:0] n_89_port_4, n_89_port_5, n_89_v;
  wire signed [`W-1:0] n_689_port_4, n_689_v;
  wire signed [`W-1:0] n_1171_port_4, n_1171_port_7, n_1171_v;
  wire signed [`W-1:0] n_127_port_3, n_127_port_6, n_127_v;
  wire signed [`W-1:0] n_259_port_5, n_259_port_8, n_259_v;
  wire signed [`W-1:0] n_1341_port_3, n_1341_port_5, n_1341_v;
  wire signed [`W-1:0] n_1072_port_5, n_1072_port_7, n_1072_v;
  wire signed [`W-1:0] n_86_port_6, n_86_port_7, n_86_v;
  wire signed [`W-1:0] n_617_port_3, n_617_port_5, n_617_v;
  wire signed [`W-1:0] n_701_port_0, n_701_port_2, n_701_port_3, n_701_port_4, n_701_v;
  wire signed [`W-1:0] n_696_port_1, n_696_port_2, n_696_port_3, n_696_port_4, n_696_v;
  wire signed [`W-1:0] n_1814_port_1, n_1814_port_2, n_1814_port_3, n_1814_v;
  wire signed [`W-1:0] reg_pcl0_port_0, reg_pcl0_port_2, reg_pcl0_port_3, reg_pcl0_v;
  wire signed [`W-1:0] n_1815_port_1, n_1815_port_2, n_1815_port_3, n_1815_v;
  wire signed [`W-1:0] reg_r0_port_0, reg_r0_port_2, reg_r0_port_3, reg_r0_v;
  wire signed [`W-1:0] n_1816_port_1, n_1816_port_2, n_1816_port_3, n_1816_v;
  wire signed [`W-1:0] reg_z0_port_0, reg_z0_port_2, reg_z0_port_3, reg_z0_v;
  wire signed [`W-1:0] n_1817_port_1, n_1817_port_2, n_1817_port_3, n_1817_v;
  wire signed [`W-1:0] reg_spl0_port_0, reg_spl0_port_2, reg_spl0_port_3, reg_spl0_v;
  wire signed [`W-1:0] n_1818_port_1, n_1818_port_2, n_1818_port_3, n_1818_v;
  wire signed [`W-1:0] reg_iyl0_port_0, reg_iyl0_port_2, reg_iyl0_port_3, reg_iyl0_v;
  wire signed [`W-1:0] n_1819_port_1, n_1819_port_2, n_1819_port_3, n_1819_v;
  wire signed [`W-1:0] reg_ixl0_port_0, reg_ixl0_port_2, reg_ixl0_port_3, reg_ixl0_v;
  wire signed [`W-1:0] n_1820_port_1, n_1820_port_2, n_1820_port_3, n_1820_v;
  wire signed [`W-1:0] reg_e0_port_0, reg_e0_port_2, reg_e0_port_3, reg_e0_v;
  wire signed [`W-1:0] n_1821_port_1, n_1821_port_2, n_1821_port_3, n_1821_v;
  wire signed [`W-1:0] reg_ee0_port_0, reg_ee0_port_2, reg_ee0_port_3, reg_ee0_v;
  wire signed [`W-1:0] n_1822_port_1, n_1822_port_2, n_1822_port_3, n_1822_v;
  wire signed [`W-1:0] reg_l0_port_0, reg_l0_port_2, reg_l0_port_3, reg_l0_v;
  wire signed [`W-1:0] n_1823_port_1, n_1823_port_2, n_1823_port_3, n_1823_v;
  wire signed [`W-1:0] reg_ll0_port_0, reg_ll0_port_2, reg_ll0_port_3, reg_ll0_v;
  wire signed [`W-1:0] n_1824_port_1, n_1824_port_2, n_1824_port_3, n_1824_v;
  wire signed [`W-1:0] reg_c0_port_0, reg_c0_port_2, reg_c0_port_3, reg_c0_v;
  wire signed [`W-1:0] n_1825_port_1, n_1825_port_2, n_1825_port_3, n_1825_v;
  wire signed [`W-1:0] reg_cc0_port_0, reg_cc0_port_2, reg_cc0_port_3, reg_cc0_v;
  wire signed [`W-1:0] n_1826_port_1, n_1826_port_2, n_1826_port_3, n_1826_v;
  wire signed [`W-1:0] reg_ff0_port_0, reg_ff0_port_2, reg_ff0_port_3, reg_ff0_v;
  wire signed [`W-1:0] n_1827_port_1, n_1827_port_2, n_1827_port_3, n_1827_v;
  wire signed [`W-1:0] reg_f0_port_0, reg_f0_port_2, reg_f0_port_3, reg_f0_v;
  wire signed [`W-1:0] n_708_port_1, n_708_port_4, n_708_port_5, n_708_port_6, n_708_port_7, n_708_port_8, n_708_port_9, n_708_port_10, n_708_port_11, n_708_port_12, n_708_port_13, n_708_port_14, n_708_port_15, n_708_port_17, n_708_v;
  wire signed [`W-1:0] n_709_port_3, n_709_port_4, n_709_port_5, n_709_v;
  wire signed [`W-1:0] n_149_port_5, n_149_port_8, n_149_v;
  wire signed [`W-1:0] n_721_port_2, n_721_port_3, n_721_port_4, n_721_v;
  wire signed [`W-1:0] n_715_port_1, n_715_port_4, n_715_port_5, n_715_port_6, n_715_port_7, n_715_port_8, n_715_port_9, n_715_port_10, n_715_port_11, n_715_port_12, n_715_port_13, n_715_port_14, n_715_port_15, n_715_port_17, n_715_v;
  wire signed [`W-1:0] n_143_port_6, n_143_port_7, n_143_v;
  wire signed [`W-1:0] reg_pcl1_port_1, reg_pcl1_port_2, reg_pcl1_port_3, reg_pcl1_v;
  wire signed [`W-1:0] n_1890_port_0, n_1890_port_2, n_1890_port_3, n_1890_v;
  wire signed [`W-1:0] reg_r1_port_1, reg_r1_port_2, reg_r1_port_3, reg_r1_v;
  wire signed [`W-1:0] n_1891_port_0, n_1891_port_2, n_1891_port_3, n_1891_v;
  wire signed [`W-1:0] reg_z1_port_1, reg_z1_port_2, reg_z1_port_3, reg_z1_v;
  wire signed [`W-1:0] n_1892_port_0, n_1892_port_2, n_1892_port_3, n_1892_v;
  wire signed [`W-1:0] reg_spl1_port_1, reg_spl1_port_2, reg_spl1_port_3, reg_spl1_v;
  wire signed [`W-1:0] n_1893_port_0, n_1893_port_2, n_1893_port_3, n_1893_v;
  wire signed [`W-1:0] reg_iyl1_port_1, reg_iyl1_port_2, reg_iyl1_port_3, reg_iyl1_v;
  wire signed [`W-1:0] n_1894_port_0, n_1894_port_2, n_1894_port_3, n_1894_v;
  wire signed [`W-1:0] reg_ixl1_port_1, reg_ixl1_port_2, reg_ixl1_port_3, reg_ixl1_v;
  wire signed [`W-1:0] n_1895_port_0, n_1895_port_2, n_1895_port_3, n_1895_v;
  wire signed [`W-1:0] reg_e1_port_1, reg_e1_port_2, reg_e1_port_3, reg_e1_v;
  wire signed [`W-1:0] n_1896_port_0, n_1896_port_2, n_1896_port_3, n_1896_v;
  wire signed [`W-1:0] reg_ee1_port_1, reg_ee1_port_2, reg_ee1_port_3, reg_ee1_v;
  wire signed [`W-1:0] n_1897_port_0, n_1897_port_2, n_1897_port_3, n_1897_v;
  wire signed [`W-1:0] reg_l1_port_1, reg_l1_port_2, reg_l1_port_3, reg_l1_v;
  wire signed [`W-1:0] n_1898_port_0, n_1898_port_2, n_1898_port_3, n_1898_v;
  wire signed [`W-1:0] reg_ll1_port_1, reg_ll1_port_2, reg_ll1_port_3, reg_ll1_v;
  wire signed [`W-1:0] n_1899_port_0, n_1899_port_2, n_1899_port_3, n_1899_v;
  wire signed [`W-1:0] reg_c1_port_1, reg_c1_port_2, reg_c1_port_3, reg_c1_v;
  wire signed [`W-1:0] n_1900_port_0, n_1900_port_2, n_1900_port_3, n_1900_v;
  wire signed [`W-1:0] reg_cc1_port_1, reg_cc1_port_2, reg_cc1_port_3, reg_cc1_v;
  wire signed [`W-1:0] n_1901_port_0, n_1901_port_2, n_1901_port_3, n_1901_v;
  wire signed [`W-1:0] reg_ff1_port_1, reg_ff1_port_2, reg_ff1_port_3, reg_ff1_v;
  wire signed [`W-1:0] n_1902_port_0, n_1902_port_2, n_1902_port_3, n_1902_v;
  wire signed [`W-1:0] reg_f1_port_1, reg_f1_port_2, reg_f1_port_3, reg_f1_v;
  wire signed [`W-1:0] n_1903_port_0, n_1903_port_2, n_1903_port_3, n_1903_v;
  wire signed [`W-1:0] n_723_port_4, n_723_v;
  wire signed [`W-1:0] n_728_port_2, n_728_port_3, n_728_port_4, n_728_v;
  wire signed [`W-1:0] n_726_port_1, n_726_port_2, n_726_port_3, n_726_port_4, n_726_port_5, n_726_v;
  wire signed [`W-1:0] n_1184_port_3, n_1184_port_4, n_1184_v;
  wire signed [`W-1:0] n_1915_port_1, n_1915_port_2, n_1915_port_3, n_1915_v;
  wire signed [`W-1:0] reg_pcl2_port_0, reg_pcl2_port_2, reg_pcl2_port_3, reg_pcl2_v;
  wire signed [`W-1:0] n_1916_port_1, n_1916_port_2, n_1916_port_3, n_1916_v;
  wire signed [`W-1:0] reg_r2_port_0, reg_r2_port_2, reg_r2_port_3, reg_r2_v;
  wire signed [`W-1:0] n_1917_port_1, n_1917_port_2, n_1917_port_3, n_1917_v;
  wire signed [`W-1:0] reg_z2_port_0, reg_z2_port_2, reg_z2_port_3, reg_z2_v;
  wire signed [`W-1:0] n_1918_port_1, n_1918_port_2, n_1918_port_3, n_1918_v;
  wire signed [`W-1:0] reg_spl2_port_0, reg_spl2_port_2, reg_spl2_port_3, reg_spl2_v;
  wire signed [`W-1:0] n_1919_port_1, n_1919_port_2, n_1919_port_3, n_1919_v;
  wire signed [`W-1:0] reg_iyl2_port_0, reg_iyl2_port_2, reg_iyl2_port_3, reg_iyl2_v;
  wire signed [`W-1:0] n_1920_port_1, n_1920_port_2, n_1920_port_3, n_1920_v;
  wire signed [`W-1:0] reg_ixl2_port_0, reg_ixl2_port_2, reg_ixl2_port_3, reg_ixl2_v;
  wire signed [`W-1:0] n_1921_port_1, n_1921_port_2, n_1921_port_3, n_1921_v;
  wire signed [`W-1:0] reg_e2_port_0, reg_e2_port_2, reg_e2_port_3, reg_e2_v;
  wire signed [`W-1:0] n_1922_port_1, n_1922_port_2, n_1922_port_3, n_1922_v;
  wire signed [`W-1:0] reg_ee2_port_0, reg_ee2_port_2, reg_ee2_port_3, reg_ee2_v;
  wire signed [`W-1:0] n_1923_port_1, n_1923_port_2, n_1923_port_3, n_1923_v;
  wire signed [`W-1:0] reg_l2_port_0, reg_l2_port_2, reg_l2_port_3, reg_l2_v;
  wire signed [`W-1:0] n_1924_port_1, n_1924_port_2, n_1924_port_3, n_1924_v;
  wire signed [`W-1:0] reg_ll2_port_0, reg_ll2_port_2, reg_ll2_port_3, reg_ll2_v;
  wire signed [`W-1:0] n_1925_port_1, n_1925_port_2, n_1925_port_3, n_1925_v;
  wire signed [`W-1:0] reg_c2_port_0, reg_c2_port_2, reg_c2_port_3, reg_c2_v;
  wire signed [`W-1:0] n_1926_port_1, n_1926_port_2, n_1926_port_3, n_1926_v;
  wire signed [`W-1:0] reg_cc2_port_0, reg_cc2_port_2, reg_cc2_port_3, reg_cc2_v;
  wire signed [`W-1:0] n_1927_port_1, n_1927_port_2, n_1927_port_3, n_1927_v;
  wire signed [`W-1:0] reg_ff2_port_0, reg_ff2_port_2, reg_ff2_port_3, reg_ff2_v;
  wire signed [`W-1:0] n_1928_port_1, n_1928_port_2, n_1928_port_3, n_1928_v;
  wire signed [`W-1:0] reg_f2_port_0, reg_f2_port_2, reg_f2_port_3, reg_f2_v;
  wire signed [`W-1:0] n_745_port_1, n_745_port_4, n_745_port_5, n_745_port_6, n_745_port_7, n_745_port_8, n_745_port_9, n_745_port_10, n_745_port_11, n_745_port_12, n_745_port_13, n_745_port_14, n_745_port_15, n_745_port_17, n_745_v;
  wire signed [`W-1:0] n_746_port_3, n_746_port_4, n_746_port_5, n_746_v;
  wire signed [`W-1:0] n_763_port_2, n_763_port_3, n_763_port_4, n_763_v;
  wire signed [`W-1:0] n_753_port_1, n_753_port_2, n_753_port_3, n_753_port_4, n_753_port_5, n_753_port_6, n_753_port_7, n_753_port_8, n_753_port_9, n_753_port_12, n_753_port_13, n_753_port_14, n_753_port_15, n_753_port_17, n_753_v;
  wire signed [`W-1:0] reg_pcl3_port_1, reg_pcl3_port_2, reg_pcl3_port_3, reg_pcl3_v;
  wire signed [`W-1:0] n_1996_port_0, n_1996_port_2, n_1996_port_3, n_1996_v;
  wire signed [`W-1:0] reg_r3_port_1, reg_r3_port_2, reg_r3_port_3, reg_r3_v;
  wire signed [`W-1:0] n_1997_port_0, n_1997_port_2, n_1997_port_3, n_1997_v;
  wire signed [`W-1:0] reg_z3_port_1, reg_z3_port_2, reg_z3_port_3, reg_z3_v;
  wire signed [`W-1:0] n_1998_port_0, n_1998_port_2, n_1998_port_3, n_1998_v;
  wire signed [`W-1:0] reg_spl3_port_1, reg_spl3_port_2, reg_spl3_port_3, reg_spl3_v;
  wire signed [`W-1:0] n_1999_port_0, n_1999_port_2, n_1999_port_3, n_1999_v;
  wire signed [`W-1:0] reg_iyl3_port_1, reg_iyl3_port_2, reg_iyl3_port_3, reg_iyl3_v;
  wire signed [`W-1:0] n_2000_port_0, n_2000_port_2, n_2000_port_3, n_2000_v;
  wire signed [`W-1:0] reg_ixl3_port_1, reg_ixl3_port_2, reg_ixl3_port_3, reg_ixl3_v;
  wire signed [`W-1:0] n_2001_port_0, n_2001_port_2, n_2001_port_3, n_2001_v;
  wire signed [`W-1:0] reg_e3_port_1, reg_e3_port_2, reg_e3_port_3, reg_e3_v;
  wire signed [`W-1:0] n_2002_port_0, n_2002_port_2, n_2002_port_3, n_2002_v;
  wire signed [`W-1:0] reg_ee3_port_1, reg_ee3_port_2, reg_ee3_port_3, reg_ee3_v;
  wire signed [`W-1:0] n_2003_port_0, n_2003_port_2, n_2003_port_3, n_2003_v;
  wire signed [`W-1:0] reg_l3_port_1, reg_l3_port_2, reg_l3_port_3, reg_l3_v;
  wire signed [`W-1:0] n_2004_port_0, n_2004_port_2, n_2004_port_3, n_2004_v;
  wire signed [`W-1:0] reg_ll3_port_1, reg_ll3_port_2, reg_ll3_port_3, reg_ll3_v;
  wire signed [`W-1:0] n_2005_port_0, n_2005_port_2, n_2005_port_3, n_2005_v;
  wire signed [`W-1:0] reg_c3_port_1, reg_c3_port_2, reg_c3_port_3, reg_c3_v;
  wire signed [`W-1:0] n_2006_port_0, n_2006_port_2, n_2006_port_3, n_2006_v;
  wire signed [`W-1:0] reg_cc3_port_1, reg_cc3_port_2, reg_cc3_port_3, reg_cc3_v;
  wire signed [`W-1:0] n_2007_port_0, n_2007_port_2, n_2007_port_3, n_2007_v;
  wire signed [`W-1:0] reg_ff3_port_1, reg_ff3_port_2, reg_ff3_port_3, reg_ff3_v;
  wire signed [`W-1:0] n_2008_port_0, n_2008_port_2, n_2008_port_3, n_2008_v;
  wire signed [`W-1:0] reg_f3_port_1, reg_f3_port_2, reg_f3_port_3, reg_f3_v;
  wire signed [`W-1:0] n_2009_port_0, n_2009_port_2, n_2009_port_3, n_2009_v;
  wire signed [`W-1:0] n_94_port_3, n_94_port_6, n_94_v;
  wire signed [`W-1:0] n_2019_port_1, n_2019_port_2, n_2019_port_3, n_2019_v;
  wire signed [`W-1:0] reg_pcl4_port_0, reg_pcl4_port_2, reg_pcl4_port_3, reg_pcl4_v;
  wire signed [`W-1:0] n_2020_port_1, n_2020_port_2, n_2020_port_3, n_2020_v;
  wire signed [`W-1:0] reg_r4_port_0, reg_r4_port_2, reg_r4_port_3, reg_r4_v;
  wire signed [`W-1:0] n_2021_port_1, n_2021_port_2, n_2021_port_3, n_2021_v;
  wire signed [`W-1:0] reg_z4_port_0, reg_z4_port_2, reg_z4_port_3, reg_z4_v;
  wire signed [`W-1:0] n_2022_port_1, n_2022_port_2, n_2022_port_3, n_2022_v;
  wire signed [`W-1:0] reg_spl4_port_0, reg_spl4_port_2, reg_spl4_port_3, reg_spl4_v;
  wire signed [`W-1:0] n_2023_port_1, n_2023_port_2, n_2023_port_3, n_2023_v;
  wire signed [`W-1:0] reg_iyl4_port_0, reg_iyl4_port_2, reg_iyl4_port_3, reg_iyl4_v;
  wire signed [`W-1:0] n_2024_port_1, n_2024_port_2, n_2024_port_3, n_2024_v;
  wire signed [`W-1:0] reg_ixl4_port_0, reg_ixl4_port_2, reg_ixl4_port_3, reg_ixl4_v;
  wire signed [`W-1:0] n_2025_port_1, n_2025_port_2, n_2025_port_3, n_2025_v;
  wire signed [`W-1:0] reg_e4_port_0, reg_e4_port_2, reg_e4_port_3, reg_e4_v;
  wire signed [`W-1:0] n_2026_port_1, n_2026_port_2, n_2026_port_3, n_2026_v;
  wire signed [`W-1:0] reg_ee4_port_0, reg_ee4_port_2, reg_ee4_port_3, reg_ee4_v;
  wire signed [`W-1:0] n_2027_port_1, n_2027_port_2, n_2027_port_3, n_2027_v;
  wire signed [`W-1:0] reg_l4_port_0, reg_l4_port_2, reg_l4_port_3, reg_l4_v;
  wire signed [`W-1:0] n_2028_port_1, n_2028_port_2, n_2028_port_3, n_2028_v;
  wire signed [`W-1:0] reg_ll4_port_0, reg_ll4_port_2, reg_ll4_port_3, reg_ll4_v;
  wire signed [`W-1:0] n_2029_port_1, n_2029_port_2, n_2029_port_3, n_2029_v;
  wire signed [`W-1:0] reg_c4_port_0, reg_c4_port_2, reg_c4_port_3, reg_c4_v;
  wire signed [`W-1:0] n_2030_port_1, n_2030_port_2, n_2030_port_3, n_2030_v;
  wire signed [`W-1:0] reg_cc4_port_0, reg_cc4_port_2, reg_cc4_port_3, reg_cc4_v;
  wire signed [`W-1:0] n_2031_port_1, n_2031_port_2, n_2031_port_3, n_2031_v;
  wire signed [`W-1:0] reg_ff4_port_0, reg_ff4_port_2, reg_ff4_port_3, reg_ff4_v;
  wire signed [`W-1:0] n_2032_port_1, n_2032_port_2, n_2032_port_3, n_2032_v;
  wire signed [`W-1:0] reg_f4_port_0, reg_f4_port_2, reg_f4_port_3, reg_f4_v;
  wire signed [`W-1:0] n_785_port_1, n_785_port_4, n_785_port_5, n_785_port_6, n_785_port_7, n_785_port_8, n_785_port_9, n_785_port_10, n_785_port_11, n_785_port_12, n_785_port_13, n_785_port_14, n_785_port_15, n_785_port_17, n_785_v;
  wire signed [`W-1:0] n_787_port_3, n_787_port_4, n_787_port_5, n_787_v;
  wire signed [`W-1:0] n_802_port_2, n_802_port_3, n_802_port_4, n_802_v;
  wire signed [`W-1:0] n_1170_port_4, n_1170_port_5, n_1170_v;
  wire signed [`W-1:0] n_799_port_1, n_799_port_4, n_799_port_5, n_799_port_6, n_799_port_7, n_799_port_8, n_799_port_9, n_799_port_10, n_799_port_11, n_799_port_12, n_799_port_13, n_799_port_14, n_799_port_15, n_799_port_17, n_799_v;
  wire signed [`W-1:0] reg_pcl5_port_1, reg_pcl5_port_2, reg_pcl5_port_3, reg_pcl5_v;
  wire signed [`W-1:0] n_2094_port_0, n_2094_port_2, n_2094_port_3, n_2094_v;
  wire signed [`W-1:0] reg_r5_port_1, reg_r5_port_2, reg_r5_port_3, reg_r5_v;
  wire signed [`W-1:0] n_2095_port_0, n_2095_port_2, n_2095_port_3, n_2095_v;
  wire signed [`W-1:0] reg_z5_port_1, reg_z5_port_2, reg_z5_port_3, reg_z5_v;
  wire signed [`W-1:0] n_2096_port_0, n_2096_port_2, n_2096_port_3, n_2096_v;
  wire signed [`W-1:0] reg_spl5_port_1, reg_spl5_port_2, reg_spl5_port_3, reg_spl5_v;
  wire signed [`W-1:0] n_2097_port_0, n_2097_port_2, n_2097_port_3, n_2097_v;
  wire signed [`W-1:0] reg_iyl5_port_1, reg_iyl5_port_2, reg_iyl5_port_3, reg_iyl5_v;
  wire signed [`W-1:0] n_2098_port_0, n_2098_port_2, n_2098_port_3, n_2098_v;
  wire signed [`W-1:0] reg_ixl5_port_1, reg_ixl5_port_2, reg_ixl5_port_3, reg_ixl5_v;
  wire signed [`W-1:0] n_2099_port_0, n_2099_port_2, n_2099_port_3, n_2099_v;
  wire signed [`W-1:0] reg_e5_port_1, reg_e5_port_2, reg_e5_port_3, reg_e5_v;
  wire signed [`W-1:0] n_2100_port_0, n_2100_port_2, n_2100_port_3, n_2100_v;
  wire signed [`W-1:0] reg_ee5_port_1, reg_ee5_port_2, reg_ee5_port_3, reg_ee5_v;
  wire signed [`W-1:0] n_2101_port_0, n_2101_port_2, n_2101_port_3, n_2101_v;
  wire signed [`W-1:0] reg_l5_port_1, reg_l5_port_2, reg_l5_port_3, reg_l5_v;
  wire signed [`W-1:0] n_2102_port_0, n_2102_port_2, n_2102_port_3, n_2102_v;
  wire signed [`W-1:0] reg_ll5_port_1, reg_ll5_port_2, reg_ll5_port_3, reg_ll5_v;
  wire signed [`W-1:0] n_2103_port_0, n_2103_port_2, n_2103_port_3, n_2103_v;
  wire signed [`W-1:0] reg_c5_port_1, reg_c5_port_2, reg_c5_port_3, reg_c5_v;
  wire signed [`W-1:0] n_2104_port_0, n_2104_port_2, n_2104_port_3, n_2104_v;
  wire signed [`W-1:0] reg_cc5_port_1, reg_cc5_port_2, reg_cc5_port_3, reg_cc5_v;
  wire signed [`W-1:0] n_2105_port_0, n_2105_port_2, n_2105_port_3, n_2105_v;
  wire signed [`W-1:0] reg_ff5_port_1, reg_ff5_port_2, reg_ff5_port_3, reg_ff5_v;
  wire signed [`W-1:0] n_2106_port_0, n_2106_port_2, n_2106_port_3, n_2106_v;
  wire signed [`W-1:0] reg_f5_port_1, reg_f5_port_2, reg_f5_port_3, reg_f5_v;
  wire signed [`W-1:0] n_2107_port_0, n_2107_port_2, n_2107_port_3, n_2107_v;
  wire signed [`W-1:0] n_2116_port_3, n_2116_v;
  wire signed [`W-1:0] n_359_port_3, n_359_port_6, n_359_v;
  wire signed [`W-1:0] n_2119_port_1, n_2119_port_2, n_2119_port_3, n_2119_v;
  wire signed [`W-1:0] reg_pcl6_port_0, reg_pcl6_port_2, reg_pcl6_port_3, reg_pcl6_v;
  wire signed [`W-1:0] n_2120_port_1, n_2120_port_2, n_2120_port_3, n_2120_v;
  wire signed [`W-1:0] reg_r6_port_0, reg_r6_port_2, reg_r6_port_3, reg_r6_v;
  wire signed [`W-1:0] n_2121_port_1, n_2121_port_2, n_2121_port_3, n_2121_v;
  wire signed [`W-1:0] reg_z6_port_0, reg_z6_port_2, reg_z6_port_3, reg_z6_v;
  wire signed [`W-1:0] n_2122_port_1, n_2122_port_2, n_2122_port_3, n_2122_v;
  wire signed [`W-1:0] reg_spl6_port_0, reg_spl6_port_2, reg_spl6_port_3, reg_spl6_v;
  wire signed [`W-1:0] n_2123_port_1, n_2123_port_2, n_2123_port_3, n_2123_v;
  wire signed [`W-1:0] reg_iyl6_port_0, reg_iyl6_port_2, reg_iyl6_port_3, reg_iyl6_v;
  wire signed [`W-1:0] n_2124_port_1, n_2124_port_2, n_2124_port_3, n_2124_v;
  wire signed [`W-1:0] reg_ixl6_port_0, reg_ixl6_port_2, reg_ixl6_port_3, reg_ixl6_v;
  wire signed [`W-1:0] n_2125_port_1, n_2125_port_2, n_2125_port_3, n_2125_v;
  wire signed [`W-1:0] reg_e6_port_0, reg_e6_port_2, reg_e6_port_3, reg_e6_v;
  wire signed [`W-1:0] n_2126_port_1, n_2126_port_2, n_2126_port_3, n_2126_v;
  wire signed [`W-1:0] reg_ee6_port_0, reg_ee6_port_2, reg_ee6_port_3, reg_ee6_v;
  wire signed [`W-1:0] n_2127_port_1, n_2127_port_2, n_2127_port_3, n_2127_v;
  wire signed [`W-1:0] reg_l6_port_0, reg_l6_port_2, reg_l6_port_3, reg_l6_v;
  wire signed [`W-1:0] n_2128_port_1, n_2128_port_2, n_2128_port_3, n_2128_v;
  wire signed [`W-1:0] reg_ll6_port_0, reg_ll6_port_2, reg_ll6_port_3, reg_ll6_v;
  wire signed [`W-1:0] n_2129_port_1, n_2129_port_2, n_2129_port_3, n_2129_v;
  wire signed [`W-1:0] reg_c6_port_0, reg_c6_port_2, reg_c6_port_3, reg_c6_v;
  wire signed [`W-1:0] n_2130_port_1, n_2130_port_2, n_2130_port_3, n_2130_v;
  wire signed [`W-1:0] reg_cc6_port_0, reg_cc6_port_2, reg_cc6_port_3, reg_cc6_v;
  wire signed [`W-1:0] n_2131_port_1, n_2131_port_2, n_2131_port_3, n_2131_v;
  wire signed [`W-1:0] reg_ff6_port_0, reg_ff6_port_2, reg_ff6_port_3, reg_ff6_v;
  wire signed [`W-1:0] n_2132_port_1, n_2132_port_2, n_2132_port_3, n_2132_v;
  wire signed [`W-1:0] reg_f6_port_0, reg_f6_port_2, reg_f6_port_3, reg_f6_v;
  wire signed [`W-1:0] n_834_port_1, n_834_port_4, n_834_port_5, n_834_port_6, n_834_port_7, n_834_port_8, n_834_port_9, n_834_port_10, n_834_port_11, n_834_port_12, n_834_port_13, n_834_port_14, n_834_port_15, n_834_port_17, n_834_v;
  wire signed [`W-1:0] n_835_port_1, n_835_port_2, n_835_port_3, n_835_v;
  wire signed [`W-1:0] n_837_port_1, n_837_port_5, n_837_port_6, n_837_port_8, n_837_port_9, n_837_v;
  wire signed [`W-1:0] n_847_port_1, n_847_port_4, n_847_port_5, n_847_port_6, n_847_port_7, n_847_port_8, n_847_port_9, n_847_port_10, n_847_port_11, n_847_port_12, n_847_port_13, n_847_port_14, n_847_port_15, n_847_port_17, n_847_v;
  wire signed [`W-1:0] n_856_port_3, n_856_port_4, n_856_port_5, n_856_v;
  wire signed [`W-1:0] reg_pcl7_port_1, reg_pcl7_port_2, reg_pcl7_port_3, reg_pcl7_v;
  wire signed [`W-1:0] n_2196_port_0, n_2196_port_2, n_2196_port_3, n_2196_v;
  wire signed [`W-1:0] reg_r7_port_1, reg_r7_port_2, reg_r7_port_3, reg_r7_v;
  wire signed [`W-1:0] n_2197_port_0, n_2197_port_2, n_2197_port_3, n_2197_v;
  wire signed [`W-1:0] reg_z7_port_1, reg_z7_port_2, reg_z7_port_3, reg_z7_v;
  wire signed [`W-1:0] n_2198_port_0, n_2198_port_2, n_2198_port_3, n_2198_v;
  wire signed [`W-1:0] reg_spl7_port_1, reg_spl7_port_2, reg_spl7_port_3, reg_spl7_v;
  wire signed [`W-1:0] n_2199_port_0, n_2199_port_2, n_2199_port_3, n_2199_v;
  wire signed [`W-1:0] reg_iyl7_port_1, reg_iyl7_port_2, reg_iyl7_port_3, reg_iyl7_v;
  wire signed [`W-1:0] n_2200_port_0, n_2200_port_2, n_2200_port_3, n_2200_v;
  wire signed [`W-1:0] reg_ixl7_port_1, reg_ixl7_port_2, reg_ixl7_port_3, reg_ixl7_v;
  wire signed [`W-1:0] n_2201_port_0, n_2201_port_2, n_2201_port_3, n_2201_v;
  wire signed [`W-1:0] reg_e7_port_1, reg_e7_port_2, reg_e7_port_3, reg_e7_v;
  wire signed [`W-1:0] n_2202_port_0, n_2202_port_2, n_2202_port_3, n_2202_v;
  wire signed [`W-1:0] reg_ee7_port_1, reg_ee7_port_2, reg_ee7_port_3, reg_ee7_v;
  wire signed [`W-1:0] n_2203_port_0, n_2203_port_2, n_2203_port_3, n_2203_v;
  wire signed [`W-1:0] reg_l7_port_1, reg_l7_port_2, reg_l7_port_3, reg_l7_v;
  wire signed [`W-1:0] n_2204_port_0, n_2204_port_2, n_2204_port_3, n_2204_v;
  wire signed [`W-1:0] reg_ll7_port_1, reg_ll7_port_2, reg_ll7_port_3, reg_ll7_v;
  wire signed [`W-1:0] n_2205_port_0, n_2205_port_2, n_2205_port_3, n_2205_v;
  wire signed [`W-1:0] reg_c7_port_1, reg_c7_port_2, reg_c7_port_3, reg_c7_v;
  wire signed [`W-1:0] n_2206_port_0, n_2206_port_2, n_2206_port_3, n_2206_v;
  wire signed [`W-1:0] reg_cc7_port_1, reg_cc7_port_2, reg_cc7_port_3, reg_cc7_v;
  wire signed [`W-1:0] n_2207_port_0, n_2207_port_2, n_2207_port_3, n_2207_v;
  wire signed [`W-1:0] reg_ff7_port_1, reg_ff7_port_2, reg_ff7_port_3, reg_ff7_v;
  wire signed [`W-1:0] n_2208_port_0, n_2208_port_2, n_2208_port_3, n_2208_v;
  wire signed [`W-1:0] reg_f7_port_1, reg_f7_port_2, reg_f7_port_3, reg_f7_v;
  wire signed [`W-1:0] n_2209_port_0, n_2209_port_2, n_2209_port_3, n_2209_v;
  wire signed [`W-1:0] n_754_port_1, n_754_port_2, n_754_port_5, n_754_v;
  wire signed [`W-1:0] n_867_port_1, n_867_port_3, n_867_port_4, n_867_port_5, n_867_v;
  wire signed [`W-1:0] n_861_port_1, n_861_port_2, n_861_port_3, n_861_v;
  wire signed [`W-1:0] n_2232_port_1, n_2232_port_2, n_2232_port_3, n_2232_v;
  wire signed [`W-1:0] reg_pch0_port_0, reg_pch0_port_2, reg_pch0_port_3, reg_pch0_v;
  wire signed [`W-1:0] n_2233_port_1, n_2233_port_2, n_2233_port_3, n_2233_v;
  wire signed [`W-1:0] reg_i0_port_0, reg_i0_port_2, reg_i0_port_3, reg_i0_v;
  wire signed [`W-1:0] n_2234_port_1, n_2234_port_2, n_2234_port_3, n_2234_v;
  wire signed [`W-1:0] reg_w0_port_0, reg_w0_port_2, reg_w0_port_3, reg_w0_v;
  wire signed [`W-1:0] n_2235_port_1, n_2235_port_2, n_2235_port_3, n_2235_v;
  wire signed [`W-1:0] reg_sph0_port_0, reg_sph0_port_2, reg_sph0_port_3, reg_sph0_v;
  wire signed [`W-1:0] n_2236_port_1, n_2236_port_2, n_2236_port_3, n_2236_v;
  wire signed [`W-1:0] reg_iyh0_port_0, reg_iyh0_port_2, reg_iyh0_port_3, reg_iyh0_v;
  wire signed [`W-1:0] n_2237_port_1, n_2237_port_2, n_2237_port_3, n_2237_v;
  wire signed [`W-1:0] reg_ixh0_port_0, reg_ixh0_port_2, reg_ixh0_port_3, reg_ixh0_v;
  wire signed [`W-1:0] n_2238_port_1, n_2238_port_2, n_2238_port_3, n_2238_v;
  wire signed [`W-1:0] reg_d0_port_0, reg_d0_port_2, reg_d0_port_3, reg_d0_v;
  wire signed [`W-1:0] n_2239_port_1, n_2239_port_2, n_2239_port_3, n_2239_v;
  wire signed [`W-1:0] reg_dd0_port_0, reg_dd0_port_2, reg_dd0_port_3, reg_dd0_v;
  wire signed [`W-1:0] n_2240_port_1, n_2240_port_2, n_2240_port_3, n_2240_v;
  wire signed [`W-1:0] reg_h0_port_0, reg_h0_port_2, reg_h0_port_3, reg_h0_v;
  wire signed [`W-1:0] n_2241_port_1, n_2241_port_2, n_2241_port_3, n_2241_v;
  wire signed [`W-1:0] reg_hh0_port_0, reg_hh0_port_2, reg_hh0_port_3, reg_hh0_v;
  wire signed [`W-1:0] n_2242_port_1, n_2242_port_2, n_2242_port_3, n_2242_v;
  wire signed [`W-1:0] reg_b0_port_0, reg_b0_port_2, reg_b0_port_3, reg_b0_v;
  wire signed [`W-1:0] n_2243_port_1, n_2243_port_2, n_2243_port_3, n_2243_v;
  wire signed [`W-1:0] reg_bb0_port_0, reg_bb0_port_2, reg_bb0_port_3, reg_bb0_v;
  wire signed [`W-1:0] n_2244_port_1, n_2244_port_2, n_2244_port_3, n_2244_v;
  wire signed [`W-1:0] reg_aa0_port_0, reg_aa0_port_2, reg_aa0_port_3, reg_aa0_v;
  wire signed [`W-1:0] n_2245_port_1, n_2245_port_2, n_2245_port_3, n_2245_v;
  wire signed [`W-1:0] reg_a0_port_0, reg_a0_port_2, reg_a0_port_3, reg_a0_v;
  wire signed [`W-1:0] n_852_port_2, n_852_port_3, n_852_port_5, n_852_port_8, n_852_port_10, n_852_v;
  wire signed [`W-1:0] n_880_port_1, n_880_port_4, n_880_port_5, n_880_port_6, n_880_port_7, n_880_port_8, n_880_port_9, n_880_port_10, n_880_port_11, n_880_port_12, n_880_port_13, n_880_port_14, n_880_port_15, n_880_port_17, n_880_v;
  wire signed [`W-1:0] n_881_port_2, n_881_port_3, n_881_port_4, n_881_v;
  wire signed [`W-1:0] n_1178_port_3, n_1178_port_6, n_1178_v;
  wire signed [`W-1:0] n_140_port_5, n_140_port_7, n_140_v;
  wire signed [`W-1:0] n_892_port_3, n_892_port_4, n_892_port_5, n_892_v;
  wire signed [`W-1:0] n_886_port_1, n_886_port_4, n_886_port_5, n_886_port_6, n_886_port_7, n_886_port_8, n_886_port_9, n_886_port_10, n_886_port_11, n_886_port_12, n_886_port_13, n_886_port_14, n_886_port_15, n_886_port_17, n_886_v;
  wire signed [`W-1:0] reg_pch1_port_1, reg_pch1_port_2, reg_pch1_port_3, reg_pch1_v;
  wire signed [`W-1:0] n_2306_port_0, n_2306_port_2, n_2306_port_3, n_2306_v;
  wire signed [`W-1:0] reg_i1_port_1, reg_i1_port_2, reg_i1_port_3, reg_i1_v;
  wire signed [`W-1:0] n_2307_port_0, n_2307_port_2, n_2307_port_3, n_2307_v;
  wire signed [`W-1:0] reg_w1_port_1, reg_w1_port_2, reg_w1_port_3, reg_w1_v;
  wire signed [`W-1:0] n_2308_port_0, n_2308_port_2, n_2308_port_3, n_2308_v;
  wire signed [`W-1:0] reg_sph1_port_1, reg_sph1_port_2, reg_sph1_port_3, reg_sph1_v;
  wire signed [`W-1:0] n_2309_port_0, n_2309_port_2, n_2309_port_3, n_2309_v;
  wire signed [`W-1:0] reg_iyh1_port_1, reg_iyh1_port_2, reg_iyh1_port_3, reg_iyh1_v;
  wire signed [`W-1:0] n_2310_port_0, n_2310_port_2, n_2310_port_3, n_2310_v;
  wire signed [`W-1:0] reg_ixh1_port_1, reg_ixh1_port_2, reg_ixh1_port_3, reg_ixh1_v;
  wire signed [`W-1:0] n_2311_port_0, n_2311_port_2, n_2311_port_3, n_2311_v;
  wire signed [`W-1:0] reg_d1_port_1, reg_d1_port_2, reg_d1_port_3, reg_d1_v;
  wire signed [`W-1:0] n_2312_port_0, n_2312_port_2, n_2312_port_3, n_2312_v;
  wire signed [`W-1:0] reg_dd1_port_1, reg_dd1_port_2, reg_dd1_port_3, reg_dd1_v;
  wire signed [`W-1:0] n_2313_port_0, n_2313_port_2, n_2313_port_3, n_2313_v;
  wire signed [`W-1:0] reg_h1_port_1, reg_h1_port_2, reg_h1_port_3, reg_h1_v;
  wire signed [`W-1:0] n_2314_port_0, n_2314_port_2, n_2314_port_3, n_2314_v;
  wire signed [`W-1:0] reg_hh1_port_1, reg_hh1_port_2, reg_hh1_port_3, reg_hh1_v;
  wire signed [`W-1:0] n_2315_port_0, n_2315_port_2, n_2315_port_3, n_2315_v;
  wire signed [`W-1:0] reg_b1_port_1, reg_b1_port_2, reg_b1_port_3, reg_b1_v;
  wire signed [`W-1:0] n_2316_port_0, n_2316_port_2, n_2316_port_3, n_2316_v;
  wire signed [`W-1:0] reg_bb1_port_1, reg_bb1_port_2, reg_bb1_port_3, reg_bb1_v;
  wire signed [`W-1:0] n_2317_port_0, n_2317_port_2, n_2317_port_3, n_2317_v;
  wire signed [`W-1:0] reg_aa1_port_1, reg_aa1_port_2, reg_aa1_port_3, reg_aa1_v;
  wire signed [`W-1:0] n_2318_port_0, n_2318_port_2, n_2318_port_3, n_2318_v;
  wire signed [`W-1:0] reg_a1_port_1, reg_a1_port_2, reg_a1_port_3, reg_a1_v;
  wire signed [`W-1:0] n_2319_port_0, n_2319_port_2, n_2319_port_3, n_2319_v;
  wire signed [`W-1:0] n_889_port_1, n_889_port_2, n_889_port_3, n_889_port_8, n_889_port_9, n_889_v;
  wire signed [`W-1:0] n_2320_port_4, n_2320_v;
  wire signed [`W-1:0] n_81_port_6, n_81_port_7, n_81_v;
  wire signed [`W-1:0] n_1076_port_5, n_1076_port_7, n_1076_v;
  wire signed [`W-1:0] n_2344_port_1, n_2344_port_2, n_2344_port_3, n_2344_v;
  wire signed [`W-1:0] reg_pch2_port_0, reg_pch2_port_2, reg_pch2_port_3, reg_pch2_v;
  wire signed [`W-1:0] n_2345_port_1, n_2345_port_2, n_2345_port_3, n_2345_v;
  wire signed [`W-1:0] reg_i2_port_0, reg_i2_port_2, reg_i2_port_3, reg_i2_v;
  wire signed [`W-1:0] n_2346_port_1, n_2346_port_2, n_2346_port_3, n_2346_v;
  wire signed [`W-1:0] reg_w2_port_0, reg_w2_port_2, reg_w2_port_3, reg_w2_v;
  wire signed [`W-1:0] n_2347_port_1, n_2347_port_2, n_2347_port_3, n_2347_v;
  wire signed [`W-1:0] reg_sph2_port_0, reg_sph2_port_2, reg_sph2_port_3, reg_sph2_v;
  wire signed [`W-1:0] n_2348_port_1, n_2348_port_2, n_2348_port_3, n_2348_v;
  wire signed [`W-1:0] reg_iyh2_port_0, reg_iyh2_port_2, reg_iyh2_port_3, reg_iyh2_v;
  wire signed [`W-1:0] n_2349_port_1, n_2349_port_2, n_2349_port_3, n_2349_v;
  wire signed [`W-1:0] reg_ixh2_port_0, reg_ixh2_port_2, reg_ixh2_port_3, reg_ixh2_v;
  wire signed [`W-1:0] n_2350_port_1, n_2350_port_2, n_2350_port_3, n_2350_v;
  wire signed [`W-1:0] reg_d2_port_0, reg_d2_port_2, reg_d2_port_3, reg_d2_v;
  wire signed [`W-1:0] n_2351_port_1, n_2351_port_2, n_2351_port_3, n_2351_v;
  wire signed [`W-1:0] reg_dd2_port_0, reg_dd2_port_2, reg_dd2_port_3, reg_dd2_v;
  wire signed [`W-1:0] n_2352_port_1, n_2352_port_2, n_2352_port_3, n_2352_v;
  wire signed [`W-1:0] reg_h2_port_0, reg_h2_port_2, reg_h2_port_3, reg_h2_v;
  wire signed [`W-1:0] n_2353_port_1, n_2353_port_2, n_2353_port_3, n_2353_v;
  wire signed [`W-1:0] reg_hh2_port_0, reg_hh2_port_2, reg_hh2_port_3, reg_hh2_v;
  wire signed [`W-1:0] n_2354_port_1, n_2354_port_2, n_2354_port_3, n_2354_v;
  wire signed [`W-1:0] reg_b2_port_0, reg_b2_port_2, reg_b2_port_3, reg_b2_v;
  wire signed [`W-1:0] n_2355_port_1, n_2355_port_2, n_2355_port_3, n_2355_v;
  wire signed [`W-1:0] reg_bb2_port_0, reg_bb2_port_2, reg_bb2_port_3, reg_bb2_v;
  wire signed [`W-1:0] n_2356_port_1, n_2356_port_2, n_2356_port_3, n_2356_v;
  wire signed [`W-1:0] reg_aa2_port_0, reg_aa2_port_2, reg_aa2_port_3, reg_aa2_v;
  wire signed [`W-1:0] n_2357_port_1, n_2357_port_2, n_2357_port_3, n_2357_v;
  wire signed [`W-1:0] reg_a2_port_0, reg_a2_port_2, reg_a2_port_3, reg_a2_v;
  wire signed [`W-1:0] n_85_port_6, n_85_port_8, n_85_v;
  wire signed [`W-1:0] n_914_port_1, n_914_port_4, n_914_port_5, n_914_port_6, n_914_port_7, n_914_port_8, n_914_port_9, n_914_port_10, n_914_port_11, n_914_port_12, n_914_port_13, n_914_port_14, n_914_port_15, n_914_port_17, n_914_v;
  wire signed [`W-1:0] n_918_port_1, n_918_port_3, n_918_port_4, n_918_port_5, n_918_v;
  wire signed [`W-1:0] n_915_port_2, n_915_port_3, n_915_port_4, n_915_v;
  wire signed [`W-1:0] n_928_port_1, n_928_port_2, n_928_port_3, n_928_v;
  wire signed [`W-1:0] n_157_port_4, n_157_port_8, n_157_v;
  wire signed [`W-1:0] n_923_port_1, n_923_port_4, n_923_port_5, n_923_port_6, n_923_port_7, n_923_port_8, n_923_port_9, n_923_port_10, n_923_port_11, n_923_port_12, n_923_port_13, n_923_port_14, n_923_port_15, n_923_port_17, n_923_v;
  wire signed [`W-1:0] reg_pch3_port_1, reg_pch3_port_2, reg_pch3_port_3, reg_pch3_v;
  wire signed [`W-1:0] n_2429_port_0, n_2429_port_2, n_2429_port_3, n_2429_v;
  wire signed [`W-1:0] reg_i3_port_1, reg_i3_port_2, reg_i3_port_3, reg_i3_v;
  wire signed [`W-1:0] n_2430_port_0, n_2430_port_2, n_2430_port_3, n_2430_v;
  wire signed [`W-1:0] reg_w3_port_1, reg_w3_port_2, reg_w3_port_3, reg_w3_v;
  wire signed [`W-1:0] n_2431_port_0, n_2431_port_2, n_2431_port_3, n_2431_v;
  wire signed [`W-1:0] reg_sph3_port_1, reg_sph3_port_2, reg_sph3_port_3, reg_sph3_v;
  wire signed [`W-1:0] n_2432_port_0, n_2432_port_2, n_2432_port_3, n_2432_v;
  wire signed [`W-1:0] reg_iyh3_port_1, reg_iyh3_port_2, reg_iyh3_port_3, reg_iyh3_v;
  wire signed [`W-1:0] n_2433_port_0, n_2433_port_2, n_2433_port_3, n_2433_v;
  wire signed [`W-1:0] reg_ixh3_port_1, reg_ixh3_port_2, reg_ixh3_port_3, reg_ixh3_v;
  wire signed [`W-1:0] n_2434_port_0, n_2434_port_2, n_2434_port_3, n_2434_v;
  wire signed [`W-1:0] reg_d3_port_1, reg_d3_port_2, reg_d3_port_3, reg_d3_v;
  wire signed [`W-1:0] n_2435_port_0, n_2435_port_2, n_2435_port_3, n_2435_v;
  wire signed [`W-1:0] reg_dd3_port_1, reg_dd3_port_2, reg_dd3_port_3, reg_dd3_v;
  wire signed [`W-1:0] n_2436_port_0, n_2436_port_2, n_2436_port_3, n_2436_v;
  wire signed [`W-1:0] reg_h3_port_1, reg_h3_port_2, reg_h3_port_3, reg_h3_v;
  wire signed [`W-1:0] n_2437_port_0, n_2437_port_2, n_2437_port_3, n_2437_v;
  wire signed [`W-1:0] reg_hh3_port_1, reg_hh3_port_2, reg_hh3_port_3, reg_hh3_v;
  wire signed [`W-1:0] n_2438_port_0, n_2438_port_2, n_2438_port_3, n_2438_v;
  wire signed [`W-1:0] reg_b3_port_1, reg_b3_port_2, reg_b3_port_3, reg_b3_v;
  wire signed [`W-1:0] n_2439_port_0, n_2439_port_2, n_2439_port_3, n_2439_v;
  wire signed [`W-1:0] reg_bb3_port_1, reg_bb3_port_2, reg_bb3_port_3, reg_bb3_v;
  wire signed [`W-1:0] n_2440_port_0, n_2440_port_2, n_2440_port_3, n_2440_v;
  wire signed [`W-1:0] reg_aa3_port_1, reg_aa3_port_2, reg_aa3_port_3, reg_aa3_v;
  wire signed [`W-1:0] n_2441_port_0, n_2441_port_2, n_2441_port_3, n_2441_v;
  wire signed [`W-1:0] reg_a3_port_1, reg_a3_port_2, reg_a3_port_3, reg_a3_v;
  wire signed [`W-1:0] n_2442_port_0, n_2442_port_2, n_2442_port_3, n_2442_v;
  wire signed [`W-1:0] n_903_port_2, n_903_port_3, n_903_port_5, n_903_port_8, n_903_port_10, n_903_v;
  wire signed [`W-1:0] n_1077_port_5, n_1077_port_8, n_1077_v;
  wire signed [`W-1:0] n_62_port_3, n_62_port_6, n_62_v;
  wire signed [`W-1:0] n_132_port_3, n_132_port_5, n_132_v;
  wire signed [`W-1:0] n_147_port_4, n_147_port_5, n_147_v;
  wire signed [`W-1:0] n_384_port_3, n_384_port_4, n_384_v;
  wire signed [`W-1:0] n_2450_port_1, n_2450_port_2, n_2450_port_3, n_2450_v;
  wire signed [`W-1:0] reg_pch4_port_0, reg_pch4_port_2, reg_pch4_port_3, reg_pch4_v;
  wire signed [`W-1:0] n_2451_port_1, n_2451_port_2, n_2451_port_3, n_2451_v;
  wire signed [`W-1:0] reg_i4_port_0, reg_i4_port_2, reg_i4_port_3, reg_i4_v;
  wire signed [`W-1:0] n_2452_port_1, n_2452_port_2, n_2452_port_3, n_2452_v;
  wire signed [`W-1:0] reg_w4_port_0, reg_w4_port_2, reg_w4_port_3, reg_w4_v;
  wire signed [`W-1:0] n_2453_port_1, n_2453_port_2, n_2453_port_3, n_2453_v;
  wire signed [`W-1:0] reg_sph4_port_0, reg_sph4_port_2, reg_sph4_port_3, reg_sph4_v;
  wire signed [`W-1:0] n_2454_port_1, n_2454_port_2, n_2454_port_3, n_2454_v;
  wire signed [`W-1:0] reg_iyh4_port_0, reg_iyh4_port_2, reg_iyh4_port_3, reg_iyh4_v;
  wire signed [`W-1:0] n_2455_port_1, n_2455_port_2, n_2455_port_3, n_2455_v;
  wire signed [`W-1:0] reg_ixh4_port_0, reg_ixh4_port_2, reg_ixh4_port_3, reg_ixh4_v;
  wire signed [`W-1:0] n_2456_port_1, n_2456_port_2, n_2456_port_3, n_2456_v;
  wire signed [`W-1:0] reg_d4_port_0, reg_d4_port_2, reg_d4_port_3, reg_d4_v;
  wire signed [`W-1:0] n_2457_port_1, n_2457_port_2, n_2457_port_3, n_2457_v;
  wire signed [`W-1:0] reg_dd4_port_0, reg_dd4_port_2, reg_dd4_port_3, reg_dd4_v;
  wire signed [`W-1:0] n_2458_port_1, n_2458_port_2, n_2458_port_3, n_2458_v;
  wire signed [`W-1:0] reg_h4_port_0, reg_h4_port_2, reg_h4_port_3, reg_h4_v;
  wire signed [`W-1:0] n_2459_port_1, n_2459_port_2, n_2459_port_3, n_2459_v;
  wire signed [`W-1:0] reg_hh4_port_0, reg_hh4_port_2, reg_hh4_port_3, reg_hh4_v;
  wire signed [`W-1:0] n_2460_port_1, n_2460_port_2, n_2460_port_3, n_2460_v;
  wire signed [`W-1:0] reg_b4_port_0, reg_b4_port_2, reg_b4_port_3, reg_b4_v;
  wire signed [`W-1:0] n_2461_port_1, n_2461_port_2, n_2461_port_3, n_2461_v;
  wire signed [`W-1:0] reg_bb4_port_0, reg_bb4_port_2, reg_bb4_port_3, reg_bb4_v;
  wire signed [`W-1:0] n_2462_port_1, n_2462_port_2, n_2462_port_3, n_2462_v;
  wire signed [`W-1:0] reg_aa4_port_0, reg_aa4_port_2, reg_aa4_port_3, reg_aa4_v;
  wire signed [`W-1:0] n_2463_port_1, n_2463_port_2, n_2463_port_3, n_2463_v;
  wire signed [`W-1:0] reg_a4_port_0, reg_a4_port_2, reg_a4_port_3, reg_a4_v;
  wire signed [`W-1:0] n_937_port_4, n_937_port_5, n_937_port_7, n_937_port_8, n_937_port_9, n_937_v;
  wire signed [`W-1:0] n_98_port_4, n_98_port_8, n_98_v;
  wire signed [`W-1:0] n_950_port_3, n_950_port_4, n_950_port_5, n_950_v;
  wire signed [`W-1:0] n_949_port_1, n_949_port_4, n_949_port_5, n_949_port_6, n_949_port_7, n_949_port_8, n_949_port_9, n_949_port_10, n_949_port_11, n_949_port_12, n_949_port_13, n_949_port_14, n_949_port_15, n_949_port_17, n_949_v;
  wire signed [`W-1:0] n_908_port_1, n_908_port_2, n_908_port_3, n_908_v;
  wire signed [`W-1:0] n_963_port_2, n_963_port_3, n_963_port_4, n_963_v;
  wire signed [`W-1:0] n_959_port_1, n_959_port_4, n_959_port_5, n_959_port_6, n_959_port_7, n_959_port_8, n_959_port_9, n_959_port_10, n_959_port_11, n_959_port_12, n_959_port_13, n_959_port_14, n_959_port_15, n_959_port_17, n_959_v;
  wire signed [`W-1:0] reg_pch5_port_1, reg_pch5_port_2, reg_pch5_port_3, reg_pch5_v;
  wire signed [`W-1:0] n_2539_port_0, n_2539_port_2, n_2539_port_3, n_2539_v;
  wire signed [`W-1:0] reg_i5_port_1, reg_i5_port_2, reg_i5_port_3, reg_i5_v;
  wire signed [`W-1:0] n_2540_port_0, n_2540_port_2, n_2540_port_3, n_2540_v;
  wire signed [`W-1:0] reg_w5_port_1, reg_w5_port_2, reg_w5_port_3, reg_w5_v;
  wire signed [`W-1:0] n_2541_port_0, n_2541_port_2, n_2541_port_3, n_2541_v;
  wire signed [`W-1:0] reg_sph5_port_1, reg_sph5_port_2, reg_sph5_port_3, reg_sph5_v;
  wire signed [`W-1:0] n_2542_port_0, n_2542_port_2, n_2542_port_3, n_2542_v;
  wire signed [`W-1:0] reg_iyh5_port_1, reg_iyh5_port_2, reg_iyh5_port_3, reg_iyh5_v;
  wire signed [`W-1:0] n_2543_port_0, n_2543_port_2, n_2543_port_3, n_2543_v;
  wire signed [`W-1:0] reg_ixh5_port_1, reg_ixh5_port_2, reg_ixh5_port_3, reg_ixh5_v;
  wire signed [`W-1:0] n_2544_port_0, n_2544_port_2, n_2544_port_3, n_2544_v;
  wire signed [`W-1:0] reg_d5_port_1, reg_d5_port_2, reg_d5_port_3, reg_d5_v;
  wire signed [`W-1:0] n_2545_port_0, n_2545_port_2, n_2545_port_3, n_2545_v;
  wire signed [`W-1:0] reg_dd5_port_1, reg_dd5_port_2, reg_dd5_port_3, reg_dd5_v;
  wire signed [`W-1:0] n_2546_port_0, n_2546_port_2, n_2546_port_3, n_2546_v;
  wire signed [`W-1:0] reg_h5_port_1, reg_h5_port_2, reg_h5_port_3, reg_h5_v;
  wire signed [`W-1:0] n_2547_port_0, n_2547_port_2, n_2547_port_3, n_2547_v;
  wire signed [`W-1:0] reg_hh5_port_1, reg_hh5_port_2, reg_hh5_port_3, reg_hh5_v;
  wire signed [`W-1:0] n_2548_port_0, n_2548_port_2, n_2548_port_3, n_2548_v;
  wire signed [`W-1:0] reg_b5_port_1, reg_b5_port_2, reg_b5_port_3, reg_b5_v;
  wire signed [`W-1:0] n_2549_port_0, n_2549_port_2, n_2549_port_3, n_2549_v;
  wire signed [`W-1:0] reg_bb5_port_1, reg_bb5_port_2, reg_bb5_port_3, reg_bb5_v;
  wire signed [`W-1:0] n_2550_port_0, n_2550_port_2, n_2550_port_3, n_2550_v;
  wire signed [`W-1:0] reg_aa5_port_1, reg_aa5_port_2, reg_aa5_port_3, reg_aa5_v;
  wire signed [`W-1:0] n_2551_port_0, n_2551_port_2, n_2551_port_3, n_2551_v;
  wire signed [`W-1:0] reg_a5_port_1, reg_a5_port_2, reg_a5_port_3, reg_a5_v;
  wire signed [`W-1:0] n_2552_port_0, n_2552_port_2, n_2552_port_3, n_2552_v;
  wire signed [`W-1:0] n_956_port_2, n_956_port_3, n_956_port_4, n_956_v;
  wire signed [`W-1:0] n_951_port_2, n_951_port_3, n_951_port_5, n_951_port_8, n_951_port_10, n_951_v;
  wire signed [`W-1:0] n_2573_port_1, n_2573_port_2, n_2573_port_3, n_2573_v;
  wire signed [`W-1:0] reg_pch6_port_0, reg_pch6_port_2, reg_pch6_port_3, reg_pch6_v;
  wire signed [`W-1:0] n_2574_port_1, n_2574_port_2, n_2574_port_3, n_2574_v;
  wire signed [`W-1:0] reg_i6_port_0, reg_i6_port_2, reg_i6_port_3, reg_i6_v;
  wire signed [`W-1:0] n_2575_port_1, n_2575_port_2, n_2575_port_3, n_2575_v;
  wire signed [`W-1:0] reg_w6_port_0, reg_w6_port_2, reg_w6_port_3, reg_w6_v;
  wire signed [`W-1:0] n_2576_port_1, n_2576_port_2, n_2576_port_3, n_2576_v;
  wire signed [`W-1:0] reg_sph6_port_0, reg_sph6_port_2, reg_sph6_port_3, reg_sph6_v;
  wire signed [`W-1:0] n_2577_port_1, n_2577_port_2, n_2577_port_3, n_2577_v;
  wire signed [`W-1:0] reg_iyh6_port_0, reg_iyh6_port_2, reg_iyh6_port_3, reg_iyh6_v;
  wire signed [`W-1:0] n_2578_port_1, n_2578_port_2, n_2578_port_3, n_2578_v;
  wire signed [`W-1:0] reg_ixh6_port_0, reg_ixh6_port_2, reg_ixh6_port_3, reg_ixh6_v;
  wire signed [`W-1:0] n_2579_port_1, n_2579_port_2, n_2579_port_3, n_2579_v;
  wire signed [`W-1:0] reg_d6_port_0, reg_d6_port_2, reg_d6_port_3, reg_d6_v;
  wire signed [`W-1:0] n_2580_port_1, n_2580_port_2, n_2580_port_3, n_2580_v;
  wire signed [`W-1:0] reg_dd6_port_0, reg_dd6_port_2, reg_dd6_port_3, reg_dd6_v;
  wire signed [`W-1:0] n_2581_port_1, n_2581_port_2, n_2581_port_3, n_2581_v;
  wire signed [`W-1:0] reg_h6_port_0, reg_h6_port_2, reg_h6_port_3, reg_h6_v;
  wire signed [`W-1:0] n_2582_port_1, n_2582_port_2, n_2582_port_3, n_2582_v;
  wire signed [`W-1:0] reg_hh6_port_0, reg_hh6_port_2, reg_hh6_port_3, reg_hh6_v;
  wire signed [`W-1:0] n_2583_port_1, n_2583_port_2, n_2583_port_3, n_2583_v;
  wire signed [`W-1:0] reg_b6_port_0, reg_b6_port_2, reg_b6_port_3, reg_b6_v;
  wire signed [`W-1:0] n_2584_port_1, n_2584_port_2, n_2584_port_3, n_2584_v;
  wire signed [`W-1:0] reg_bb6_port_0, reg_bb6_port_2, reg_bb6_port_3, reg_bb6_v;
  wire signed [`W-1:0] n_2585_port_1, n_2585_port_2, n_2585_port_3, n_2585_v;
  wire signed [`W-1:0] reg_aa6_port_0, reg_aa6_port_2, reg_aa6_port_3, reg_aa6_v;
  wire signed [`W-1:0] n_2586_port_1, n_2586_port_2, n_2586_port_3, n_2586_v;
  wire signed [`W-1:0] reg_a6_port_0, reg_a6_port_2, reg_a6_port_3, reg_a6_v;
  wire signed [`W-1:0] _reset_port_1, _reset_v;
  wire signed [`W-1:0] n_980_port_1, n_980_port_4, n_980_port_5, n_980_port_6, n_980_port_7, n_980_port_8, n_980_port_9, n_980_port_10, n_980_port_11, n_980_port_12, n_980_port_13, n_980_port_14, n_980_port_15, n_980_port_17, n_980_v;
  wire signed [`W-1:0] n_981_port_1, n_981_port_2, n_981_port_3, n_981_v;
  wire signed [`W-1:0] n_2617_port_4, n_2617_v;
  wire signed [`W-1:0] n_985_port_1, n_985_port_4, n_985_port_5, n_985_port_6, n_985_port_7, n_985_port_8, n_985_port_9, n_985_port_10, n_985_port_11, n_985_port_12, n_985_port_13, n_985_port_14, n_985_port_15, n_985_port_17, n_985_v;
  wire signed [`W-1:0] n_983_port_4, n_983_port_5, n_983_port_7, n_983_port_8, n_983_port_9, n_983_v;
  wire signed [`W-1:0] reg_pch7_port_1, reg_pch7_port_2, reg_pch7_port_3, reg_pch7_v;
  wire signed [`W-1:0] n_2643_port_0, n_2643_port_2, n_2643_port_3, n_2643_v;
  wire signed [`W-1:0] reg_i7_port_1, reg_i7_port_2, reg_i7_port_3, reg_i7_v;
  wire signed [`W-1:0] n_2644_port_0, n_2644_port_2, n_2644_port_3, n_2644_v;
  wire signed [`W-1:0] reg_w7_port_1, reg_w7_port_2, reg_w7_port_3, reg_w7_v;
  wire signed [`W-1:0] n_2645_port_0, n_2645_port_2, n_2645_port_3, n_2645_v;
  wire signed [`W-1:0] reg_sph7_port_1, reg_sph7_port_2, reg_sph7_port_3, reg_sph7_v;
  wire signed [`W-1:0] n_2646_port_0, n_2646_port_2, n_2646_port_3, n_2646_v;
  wire signed [`W-1:0] reg_iyh7_port_1, reg_iyh7_port_2, reg_iyh7_port_3, reg_iyh7_v;
  wire signed [`W-1:0] n_2647_port_0, n_2647_port_2, n_2647_port_3, n_2647_v;
  wire signed [`W-1:0] reg_ixh7_port_1, reg_ixh7_port_2, reg_ixh7_port_3, reg_ixh7_v;
  wire signed [`W-1:0] n_2648_port_0, n_2648_port_2, n_2648_port_3, n_2648_v;
  wire signed [`W-1:0] reg_d7_port_1, reg_d7_port_2, reg_d7_port_3, reg_d7_v;
  wire signed [`W-1:0] n_2649_port_0, n_2649_port_2, n_2649_port_3, n_2649_v;
  wire signed [`W-1:0] reg_dd7_port_1, reg_dd7_port_2, reg_dd7_port_3, reg_dd7_v;
  wire signed [`W-1:0] n_2650_port_0, n_2650_port_2, n_2650_port_3, n_2650_v;
  wire signed [`W-1:0] reg_h7_port_1, reg_h7_port_2, reg_h7_port_3, reg_h7_v;
  wire signed [`W-1:0] n_2651_port_0, n_2651_port_2, n_2651_port_3, n_2651_v;
  wire signed [`W-1:0] reg_hh7_port_1, reg_hh7_port_2, reg_hh7_port_3, reg_hh7_v;
  wire signed [`W-1:0] n_2652_port_0, n_2652_port_2, n_2652_port_3, n_2652_v;
  wire signed [`W-1:0] reg_b7_port_1, reg_b7_port_2, reg_b7_port_3, reg_b7_v;
  wire signed [`W-1:0] n_2653_port_0, n_2653_port_2, n_2653_port_3, n_2653_v;
  wire signed [`W-1:0] reg_bb7_port_1, reg_bb7_port_2, reg_bb7_port_3, reg_bb7_v;
  wire signed [`W-1:0] n_2654_port_0, n_2654_port_2, n_2654_port_3, n_2654_v;
  wire signed [`W-1:0] reg_aa7_port_1, reg_aa7_port_2, reg_aa7_port_3, reg_aa7_v;
  wire signed [`W-1:0] n_2655_port_0, n_2655_port_2, n_2655_port_3, n_2655_v;
  wire signed [`W-1:0] reg_a7_port_1, reg_a7_port_2, reg_a7_port_3, reg_a7_v;
  wire signed [`W-1:0] n_2656_port_0, n_2656_port_2, n_2656_port_3, n_2656_v;
  wire signed [`W-1:0] n_988_port_1, n_988_port_2, n_988_port_4, n_988_port_5, n_988_v;
  wire signed [`W-1:0] n_1001_port_2, n_1001_port_3, n_1001_port_4, n_1001_v;
  wire signed [`W-1:0] n_995_port_2, n_995_port_3, n_995_port_4, n_995_port_8, n_995_port_10, n_995_v;
  wire signed [`W-1:0] n_1009_port_4, n_1009_v;
  wire signed [`W-1:0] n_408_port_4, n_408_port_6, n_408_v;
  wire signed [`W-1:0] n_2700_port_4, n_2700_v;
  wire signed [`W-1:0] n_2701_port_4, n_2701_v;
  wire signed [`W-1:0] n_2702_port_4, n_2702_v;
  wire signed [`W-1:0] n_2703_port_4, n_2703_v;
  wire signed [`W-1:0] n_2704_port_4, n_2704_v;
  wire signed [`W-1:0] n_2705_port_4, n_2705_v;
  wire signed [`W-1:0] n_1014_port_4, n_1014_v;
  wire signed [`W-1:0] n_1017_port_4, n_1017_v;
  wire signed [`W-1:0] n_1018_port_4, n_1018_v;
  wire signed [`W-1:0] n_1020_port_4, n_1020_v;
  wire signed [`W-1:0] n_118_port_4, n_118_port_7, n_118_v;
  wire signed [`W-1:0] n_169_port_3, n_169_port_6, n_169_v;
  wire signed [`W-1:0] n_1204_port_3, n_1204_port_5, n_1204_v;
  wire signed [`W-1:0] n_902_port_0, n_902_port_1, n_902_port_2, n_902_port_3, n_902_port_4, n_902_port_5, n_902_port_6, n_902_port_7, n_902_port_8, n_902_port_9, n_902_port_10, n_902_port_11, n_902_port_13, n_902_port_15, n_902_v;
  wire signed [`W-1:0] n_769_port_1, n_769_port_2, n_769_port_3, n_769_v;
  wire signed [`W-1:0] n_906_port_0, n_906_port_1, n_906_port_2, n_906_port_3, n_906_port_4, n_906_port_5, n_906_port_6, n_906_port_7, n_906_port_8, n_906_port_9, n_906_port_10, n_906_port_11, n_906_port_13, n_906_port_15, n_906_v;
  wire signed [`W-1:0] n_1217_port_2, n_1217_port_4, n_1217_v;
  wire signed [`W-1:0] n_913_port_0, n_913_port_1, n_913_port_3, n_913_v;
  wire signed [`W-1:0] n_328_port_2, n_328_port_3, n_328_v;
  wire signed [`W-1:0] n_775_port_1, n_775_port_3, n_775_port_4, n_775_port_5, n_775_port_6, n_775_port_7, n_775_port_8, n_775_port_9, n_775_port_10, n_775_port_11, n_775_port_12, n_775_port_13, n_775_port_14, n_775_port_15, n_775_v;
  wire signed [`W-1:0] n_1061_v;
  wire signed [`W-1:0] n_2775_port_0, n_2775_v;
  wire signed [`W-1:0] n_2776_port_0, n_2776_v;
  wire signed [`W-1:0] n_225_port_2, n_225_port_3, n_225_v;
  wire signed [`W-1:0] n_475_port_7, n_475_v;
  wire signed [`W-1:0] n_776_port_0, n_776_port_1, n_776_port_2, n_776_port_3, n_776_port_4, n_776_port_5, n_776_port_6, n_776_port_7, n_776_port_8, n_776_port_9, n_776_port_10, n_776_port_11, n_776_port_13, n_776_port_15, n_776_v;
  wire signed [`W-1:0] n_1383_port_2, n_1383_port_4, n_1383_v;
  wire signed [`W-1:0] n_784_port_0, n_784_port_1, n_784_port_3, n_784_v;
  wire signed [`W-1:0] n_1090_port_2, n_1090_port_4, n_1090_v;
  wire signed [`W-1:0] n_929_port_1, n_929_port_2, n_929_port_3, n_929_v;
  wire signed [`W-1:0] n_541_port_2, n_541_port_3, n_541_v;
  wire signed [`W-1:0] n_1405_port_2, n_1405_port_3, n_1405_v;
  wire signed [`W-1:0] n_1327_port_2, n_1327_port_3, n_1327_v;
  wire signed [`W-1:0] n_934_port_1, n_934_port_3, n_934_port_4, n_934_port_5, n_934_port_6, n_934_port_7, n_934_port_8, n_934_port_9, n_934_port_10, n_934_port_11, n_934_port_12, n_934_port_13, n_934_port_14, n_934_port_15, n_934_v;
  wire signed [`W-1:0] n_1098_port_2, n_1098_port_4, n_1098_v;
  wire signed [`W-1:0] n_935_port_0, n_935_port_1, n_935_port_2, n_935_port_3, n_935_port_4, n_935_port_5, n_935_port_6, n_935_port_7, n_935_port_8, n_935_port_9, n_935_port_10, n_935_port_11, n_935_port_13, n_935_port_15, n_935_v;
  wire signed [`W-1:0] n_161_port_2, n_161_port_4, n_161_v;
  wire signed [`W-1:0] n_948_port_0, n_948_port_1, n_948_port_3, n_948_v;
  wire signed [`W-1:0] n_146_port_2, n_146_port_4, n_146_v;
  wire signed [`W-1:0] n_700_port_1, n_700_port_2, n_700_port_3, n_700_v;
  wire signed [`W-1:0] n_804_port_1, n_804_port_2, n_804_port_3, n_804_v;
  wire signed [`W-1:0] n_702_port_0, n_702_port_1, n_702_port_2, n_702_port_3, n_702_port_4, n_702_port_5, n_702_port_6, n_702_port_7, n_702_port_8, n_702_port_9, n_702_port_10, n_702_port_11, n_702_port_13, n_702_port_15, n_702_v;
  wire signed [`W-1:0] n_807_port_1, n_807_port_3, n_807_port_4, n_807_port_5, n_807_port_6, n_807_port_7, n_807_port_8, n_807_port_9, n_807_port_10, n_807_port_11, n_807_port_12, n_807_port_13, n_807_port_14, n_807_port_15, n_807_v;
  wire signed [`W-1:0] n_964_port_1, n_964_port_2, n_964_port_3, n_964_v;
  wire signed [`W-1:0] n_707_port_0, n_707_port_1, n_707_port_3, n_707_v;
  wire signed [`W-1:0] n_809_port_0, n_809_port_1, n_809_port_2, n_809_port_3, n_809_port_4, n_809_port_5, n_809_port_6, n_809_port_7, n_809_port_8, n_809_port_9, n_809_port_10, n_809_port_11, n_809_port_13, n_809_port_15, n_809_v;
  wire signed [`W-1:0] n_833_port_0, n_833_port_1, n_833_port_3, n_833_v;
  wire signed [`W-1:0] n_970_port_1, n_970_port_3, n_970_port_4, n_970_port_5, n_970_port_6, n_970_port_7, n_970_port_8, n_970_port_9, n_970_port_10, n_970_port_11, n_970_port_12, n_970_port_13, n_970_port_14, n_970_port_15, n_970_v;
  wire signed [`W-1:0] n_973_port_0, n_973_port_1, n_973_port_2, n_973_port_3, n_973_port_4, n_973_port_5, n_973_port_6, n_973_port_7, n_973_port_8, n_973_port_9, n_973_port_10, n_973_port_11, n_973_port_13, n_973_port_15, n_973_v;
  wire signed [`W-1:0] n_979_port_0, n_979_port_1, n_979_port_3, n_979_v;
  wire signed [`W-1:0] n_857_port_1, n_857_port_2, n_857_port_3, n_857_v;
  wire signed [`W-1:0] n_1649_port_2, n_1649_port_4, n_1649_v;
  wire signed [`W-1:0] n_722_port_1, n_722_port_2, n_722_port_3, n_722_v;
  wire signed [`W-1:0] n_994_port_1, n_994_port_2, n_994_port_3, n_994_v;
  wire signed [`W-1:0] n_864_port_1, n_864_port_3, n_864_port_4, n_864_port_5, n_864_port_6, n_864_port_7, n_864_port_8, n_864_port_9, n_864_port_10, n_864_port_11, n_864_port_12, n_864_port_13, n_864_port_14, n_864_port_15, n_864_v;
  wire signed [`W-1:0] n_732_port_1, n_732_port_3, n_732_port_4, n_732_port_5, n_732_port_6, n_732_port_7, n_732_port_8, n_732_port_9, n_732_port_10, n_732_port_11, n_732_port_12, n_732_port_13, n_732_port_14, n_732_port_15, n_732_v;
  wire signed [`W-1:0] n_999_port_1, n_999_port_3, n_999_port_4, n_999_port_5, n_999_port_6, n_999_port_7, n_999_port_8, n_999_port_9, n_999_port_10, n_999_port_11, n_999_port_12, n_999_port_13, n_999_port_14, n_999_port_15, n_999_v;
  wire signed [`W-1:0] n_870_port_0, n_870_port_1, n_870_port_2, n_870_port_3, n_870_port_4, n_870_port_5, n_870_port_6, n_870_port_7, n_870_port_8, n_870_port_9, n_870_port_10, n_870_port_11, n_870_port_13, n_870_port_15, n_870_v;
  wire signed [`W-1:0] n_738_port_0, n_738_port_1, n_738_port_2, n_738_port_3, n_738_port_4, n_738_port_5, n_738_port_6, n_738_port_7, n_738_port_8, n_738_port_9, n_738_port_10, n_738_port_11, n_738_port_13, n_738_port_15, n_738_v;
  wire signed [`W-1:0] n_879_port_0, n_879_port_1, n_879_port_3, n_879_v;
  wire signed [`W-1:0] n_1044_port_2, n_1044_port_3, n_1044_v;
  wire signed [`W-1:0] n_744_port_0, n_744_port_1, n_744_port_3, n_744_v;
  wire signed [`W-1:0] n_893_port_1, n_893_port_2, n_893_port_3, n_893_v;

  wire n_2041_v;
  wire n_2037_v;
  wire n_792_v;
  wire n_1069_v;
  wire n_1042_v;
  wire n_1039_v;
  wire _rd_v;
  wire n_1249_v;
  wire n_95_v;
  wire n_1346_v;
  wire n_371_v;
  wire n_781_v;
  wire n_3421_v;
  wire n_2036_v;
  wire n_3420_v;
  wire n_608_v;
  wire n_220_v;
  wire n_706_v;
  wire n_3366_v;
  wire n_911_v;
  wire n_3493_v;
  wire n_823_v;
  wire n_794_v;
  wire n_909_v;
  wire n_3494_v;
  wire n_704_v;
  wire n_3367_v;
  wire n_170_v;
  wire n_1241_v;
  wire m4_v;
  wire n_1359_v;
  wire n_1358_v;
  wire n_100_v;
  wire _mreq_v;
  wire n_383_v;
  wire n_1362_v;
  wire n_2937_v;
  wire n_373_v;
  wire n_375_v;
  wire n_1156_v;
  wire n_99_v;
  wire n_2367_v;
  wire n_250_v;
  wire n_1309_v;
  wire n_254_v;
  wire n_1505_v;
  wire n_588_v;
  wire n_1834_v;
  wire n_3372_v;
  wire n_1507_v;
  wire n_2364_v;
  wire n_2396_v;
  wire n_1838_v;
  wire n_795_v;
  wire n_705_v;
  wire n_3375_v;
  wire n_800_v;
  wire n_3424_v;
  wire n_910_v;
  wire n_3499_v;
  wire n_2363_v;
  wire n_3498_v;
  wire n_1833_v;
  wire n_3374_v;
  wire n_1247_v;
  wire m5_v;
  wire n_1312_v;
  wire n_192_v;
  wire n_1644_v;
  wire n_600_v;
  wire n_1651_v;
  wire n_602_v;
  wire n_1510_v;
  wire n_1365_v;
  wire n_1364_v;
  wire n_1511_v;
  wire n_465_v;
  wire n_2084_v;
  wire n_3415_v;
  wire n_1318_v;
  wire n_177_v;
  wire n_829_v;
  wire n_3412_v;
  wire n_2061_v;
  wire n_3416_v;
  wire n_3411_v;
  wire n_2087_v;
  wire n_3426_v;
  wire n_2063_v;
  wire n_3407_v;
  wire n_2086_v;
  wire n_797_v;
  wire n_2066_v;
  wire n_3414_v;
  wire n_2386_v;
  wire n_2421_v;
  wire n_2091_v;
  wire ab2_v;
  wire n_1514_v;
  wire n_589_v;
  wire n_924_v;
  wire n_925_v;
  wire n_2388_v;
  wire n_3509_v;
  wire n_376_v;
  wire n_378_v;
  wire n_2064_v;
  wire n_3413_v;
  wire n_3409_v;
  wire n_1658_v;
  wire n_1674_v;
  wire n_2390_v;
  wire n_3511_v;
  wire n_2108_v;
  wire n_926_v;
  wire n_3506_v;
  wire n_2062_v;
  wire n_3408_v;
  wire n_1317_v;
  wire n_267_v;
  wire n_1661_v;
  wire n_750_v;
  wire n_788_v;
  wire n_3428_v;
  wire n_1408_v;
  wire n_2971_v;
  wire n_1665_v;
  wire n_627_v;
  wire n_2109_v;
  wire n_822_v;
  wire n_2111_v;
  wire n_821_v;
  wire n_1316_v;
  wire n_263_v;
  wire n_1369_v;
  wire n_1368_v;
  wire n_2112_v;
  wire n_820_v;
  wire n_1202_v;
  wire n_133_v;
  wire n_2420_v;
  wire n_3508_v;
  wire n_2419_v;
  wire n_921_v;
  wire n_2393_v;
  wire n_2330_v;
  wire n_2398_v;
  wire n_3513_v;
  wire n_379_v;
  wire n_1371_v;
  wire n_2395_v;
  wire n_805_v;
  wire n_3429_v;
  wire n_2397_v;
  wire n_1679_v;
  wire n_603_v;
  wire n_2444_v;
  wire n_801_v;
  wire n_3430_v;
  wire n_2110_v;
  wire n_831_v;
  wire n_1418_v;
  wire n_436_v;
  wire n_832_v;
  wire n_920_v;
  wire n_2426_v;
  wire n_896_v;
  wire n_2115_v;
  wire n_824_v;
  wire n_1680_v;
  wire n_604_v;
  wire n_718_v;
  wire n_3381_v;
  wire n_733_v;
  wire n_931_v;
  wire n_3514_v;
  wire n_927_v;
  wire n_3515_v;
  wire ab3_v;
  wire n_1374_v;
  wire n_1373_v;
  wire n_1270_v;
  wire n_103_v;
  wire n_1372_v;
  wire _m1_v;
  wire n_386_v;
  wire n_107_v;
  wire n_382_v;
  wire n_1377_v;
  wire n_1056_v;
  wire n_59_v;
  wire n_1328_v;
  wire n_126_v;
  wire n_2117_v;
  wire n_1379_v;
  wire n_1885_v;
  wire n_3385_v;
  wire n_1883_v;
  wire n_3383_v;
  wire n_1154_v;
  wire _t1_v;
  wire n_1035_v;
  wire _halt_v;
  wire m6_v;
  wire n_1378_v;
  wire n_1376_v;
  wire n_1045_v;
  wire n_64_v;
  wire n_388_v;
  wire n_385_v;
  wire n_106_v;
  wire n_1905_v;
  wire n_815_v;
  wire n_3432_v;
  wire n_941_v;
  wire n_3518_v;
  wire n_812_v;
  wire n_3433_v;
  wire n_938_v;
  wire n_3519_v;
  wire n_1533_v;
  wire n_502_v;
  wire n_1181_v;
  wire n_2820_v;
  wire n_1707_v;
  wire n_1381_v;
  wire n_393_v;
  wire n_1047_v;
  wire n_54_v;
  wire n_1387_v;
  wire n_247_v;
  wire n_725_v;
  wire n_3389_v;
  wire n_2471_v;
  wire n_2445_v;
  wire n_3522_v;
  wire n_1074_v;
  wire n_1038_v;
  wire n_2140_v;
  wire n_2468_v;
  wire n_954_v;
  wire n_2491_v;
  wire n_719_v;
  wire n_3390_v;
  wire n_1884_v;
  wire n_1912_v;
  wire n_2137_v;
  wire n_2160_v;
  wire n_2499_v;
  wire n_3521_v;
  wire n_2498_v;
  wire n_3523_v;
  wire n_939_v;
  wire n_3529_v;
  wire n_2500_v;
  wire n_2494_v;
  wire n_2467_v;
  wire n_3527_v;
  wire n_392_v;
  wire n_1386_v;
  wire n_2506_v;
  wire n_2492_v;
  wire n_1428_v;
  wire n_452_v;
  wire n_814_v;
  wire n_3436_v;
  wire n_2509_v;
  wire n_3525_v;
  wire n_2136_v;
  wire n_3435_v;
  wire ab1_v;
  wire n_1330_v;
  wire n_1075_v;
  wire n_87_v;
  wire n_1394_v;
  wire n_1390_v;
  wire n_1086_v;
  wire n_83_v;
  wire n_1440_v;
  wire _rfsh_v;
  wire n_1186_v;
  wire n_101_v;
  wire n_1088_v;
  wire n_1036_v;
  wire n_1717_v;
  wire n_1071_v;
  wire n_90_v;
  wire n_1434_v;
  wire n_456_v;
  wire n_1430_v;
  wire n_1913_v;
  wire n_1753_v;
  wire n_961_v;
  wire n_3534_v;
  wire n_1117_v;
  wire n_1058_v;
  wire n_1280_v;
  wire n_228_v;
  wire n_2181_v;
  wire n_1216_v;
  wire _t3_v;
  wire n_851_v;
  wire n_3441_v;
  wire n_1441_v;
  wire n_1439_v;
  wire n_1288_v;
  wire n_2882_v;
  wire _wr_v;
  wire n_1118_v;
  wire n_108_v;
  wire n_1203_v;
  wire n_1455_v;
  wire n_395_v;
  wire n_2533_v;
  wire n_3536_v;
  wire n_1286_v;
  wire n_204_v;
  wire n_743_v;
  wire n_3392_v;
  wire n_2532_v;
  wire n_957_v;
  wire n_2185_v;
  wire n_3443_v;
  wire n_2182_v;
  wire n_2163_v;
  wire n_2189_v;
  wire n_3440_v;
  wire n_741_v;
  wire n_3393_v;
  wire n_2191_v;
  wire n_2184_v;
  wire n_1932_v;
  wire n_734_v;
  wire n_1113_v;
  wire n_119_v;
  wire n_2555_v;
  wire n_2210_v;
  wire n_3439_v;
  wire n_1120_v;
  wire n_122_v;
  wire n_1748_v;
  wire ab0_v;
  wire n_2215_v;
  wire n_2217_v;
  wire n_3444_v;
  wire n_2214_v;
  wire n_2158_v;
  wire n_1295_v;
  wire _t4_v;
  wire n_965_v;
  wire n_3541_v;
  wire _busak_v;
  wire n_1214_v;
  wire n_142_v;
  wire n_2553_v;
  wire n_2569_v;
  wire n_962_v;
  wire n_3542_v;
  wire n_972_v;
  wire n_767_v;
  wire n_1065_v;
  wire n_69_v;
  wire n_1933_v;
  wire n_747_v;
  wire n_2554_v;
  wire n_3546_v;
  wire n_1193_v;
  wire n_188_v;
  wire n_859_v;
  wire n_1209_v;
  wire m2_v;
  wire n_1451_v;
  wire n_607_v;
  wire n_1936_v;
  wire n_1968_v;
  wire n_858_v;
  wire n_3452_v;
  wire n_1940_v;
  wire n_853_v;
  wire n_3453_v;
  wire n_1736_v;
  wire n_1785_v;
  wire n_1961_v;
  wire n_735_v;
  wire n_1579_v;
  wire n_575_v;
  wire n_2556_v;
  wire n_3547_v;
  wire n_1063_v;
  wire n_978_v;
  wire n_1962_v;
  wire n_757_v;
  wire n_2560_v;
  wire n_2496_v;
  wire n_2564_v;
  wire n_3551_v;
  wire n_1762_v;
  wire n_1119_v;
  wire n_131_v;
  wire n_1064_v;
  wire n_1037_v;
  wire n_1471_v;
  wire n_1462_v;
  wire n_1964_v;
  wire n_740_v;
  wire n_742_v;
  wire n_3396_v;
  wire n_1737_v;
  wire n_680_v;
  wire n_1935_v;
  wire n_3395_v;
  wire n_1130_v;
  wire n_111_v;
  wire n_1194_v;
  wire _t5_v;
  wire n_1593_v;
  wire n_651_v;
  wire n_1766_v;
  wire n_643_v;
  wire n_977_v;
  wire n_3549_v;
  wire n_2565_v;
  wire n_817_v;
  wire n_2561_v;
  wire n_1292_v;
  wire n_110_v;
  wire n_975_v;
  wire n_3550_v;
  wire n_2563_v;
  wire n_1097_v;
  wire n_93_v;
  wire n_1473_v;
  wire n_232_v;
  wire n_1769_v;
  wire n_646_v;
  wire n_1335_v;
  wire n_162_v;
  wire n_2568_v;
  wire n_2229_v;
  wire n_1191_v;
  wire _t6_v;
  wire n_2594_v;
  wire n_968_v;
  wire n_2571_v;
  wire n_943_v;
  wire n_1093_v;
  wire n_105_v;
  wire n_1094_v;
  wire n_66_v;
  wire n_2591_v;
  wire n_1003_v;
  wire n_1103_v;
  wire n_1040_v;
  wire n_1223_v;
  wire n_165_v;
  wire n_1751_v;
  wire n_976_v;
  wire n_3554_v;
  wire n_2590_v;
  wire n_3553_v;
  wire n_1068_v;
  wire n_80_v;
  wire n_1226_v;
  wire n_1207_v;
  wire n_1779_v;
  wire n_641_v;
  wire n_1965_v;
  wire n_1969_v;
  wire n_1966_v;
  wire n_877_v;
  wire n_3463_v;
  wire n_875_v;
  wire n_878_v;
  wire n_1788_v;
  wire n_693_v;
  wire n_873_v;
  wire n_3464_v;
  wire n_2224_v;
  wire n_3467_v;
  wire _iorq_v;
  wire n_1599_v;
  wire n_194_v;
  wire n_2616_v;
  wire ab4_v;
  wire n_760_v;
  wire n_3399_v;
  wire n_987_v;
  wire n_3558_v;
  wire n_1242_v;
  wire n_1104_v;
  wire n_1790_v;
  wire n_684_v;
  wire n_1301_v;
  wire n_222_v;
  wire n_2226_v;
  wire n_3469_v;
  wire n_679_v;
  wire n_678_v;
  wire n_1786_v;
  wire n_692_v;
  wire n_2254_v;
  wire n_2230_v;
  wire n_2186_v;
  wire n_1607_v;
  wire n_590_v;
  wire n_2613_v;
  wire n_2615_v;
  wire n_2637_v;
  wire n_3560_v;
  wire n_2636_v;
  wire n_653_v;
  wire n_652_v;
  wire n_2641_v;
  wire n_1620_v;
  wire n_574_v;
  wire n_2251_v;
  wire n_2279_v;
  wire n_2227_v;
  wire n_3471_v;
  wire n_1991_v;
  wire n_3401_v;
  wire n_2665_v;
  wire n_2663_v;
  wire n_3557_v;
  wire n_2231_v;
  wire n_2662_v;
  wire n_3562_v;
  wire n_2664_v;
  wire n_2658_v;
  wire n_2247_v;
  wire n_1990_v;
  wire n_1970_v;
  wire n_1989_v;
  wire n_3404_v;
  wire n_1617_v;
  wire n_618_v;
  wire n_2639_v;
  wire n_1004_v;
  wire n_1392_v;
  wire n_65_v;
  wire n_874_v;
  wire n_3473_v;
  wire n_2673_v;
  wire n_3564_v;
  wire n_2250_v;
  wire n_3472_v;
  wire n_996_v;
  wire n_3569_v;
  wire n_990_v;
  wire n_3570_v;
  wire n_868_v;
  wire n_2273_v;
  wire n_844_v;
  wire n_1625_v;
  wire n_552_v;
  wire n_2010_v;
  wire n_655_v;
  wire n_654_v;
  wire n_1243_v;
  wire n_397_v;
  wire n_1393_v;
  wire n_656_v;
  wire n_657_v;
  wire n_659_v;
  wire n_658_v;
  wire n_1245_v;
  wire n_1338_v;
  wire n_1336_v;
  wire n_660_v;
  wire n_661_v;
  wire n_663_v;
  wire n_662_v;
  wire n_1482_v;
  wire n_479_v;
  wire n_1340_v;
  wire n_326_v;
  wire n_664_v;
  wire n_665_v;
  wire n_771_v;
  wire n_3405_v;
  wire n_761_v;
  wire n_3406_v;
  wire n_667_v;
  wire n_666_v;
  wire n_1344_v;
  wire m1_v;
  wire n_1631_v;
  wire n_553_v;
  wire n_888_v;
  wire n_3477_v;
  wire n_668_v;
  wire n_669_v;
  wire n_671_v;
  wire n_670_v;
  wire n_1401_v;
  wire n_1385_v;
  wire n_1149_v;
  wire n_129_v;
  wire n_672_v;
  wire n_673_v;
  wire n_675_v;
  wire n_674_v;
  wire n_1638_v;
  wire n_612_v;
  wire n_1627_v;
  wire n_558_v;
  wire n_676_v;
  wire n_677_v;
  wire n_1339_v;
  wire n_327_v;
  wire n_1008_v;
  wire n_827_v;
  wire n_2680_v;
  wire n_3581_v;
  wire n_1070_v;
  wire n_78_v;
  wire n_1492_v;
  wire n_548_v;
  wire n_2685_v;
  wire n_2677_v;
  wire n_3579_v;
  wire n_1634_v;
  wire n_551_v;
  wire n_2682_v;
  wire n_3583_v;
  wire n_1804_v;
  wire n_2300_v;
  wire n_3479_v;
  wire n_2683_v;
  wire n_2659_v;
  wire n_2299_v;
  wire n_2280_v;
  wire n_1626_v;
  wire n_549_v;
  wire n_2687_v;
  wire n_3584_v;
  wire n_2688_v;
  wire n_830_v;
  wire n_2686_v;
  wire n_2014_v;
  wire n_2044_v;
  wire n_1400_v;
  wire n_1354_v;
  wire n_1007_v;
  wire n_2693_v;
  wire n_989_v;
  wire n_2696_v;
  wire n_2695_v;
  wire n_1801_v;
  wire n_1303_v;
  wire n_265_v;
  wire n_2321_v;
  wire n_2699_v;
  wire n_883_v;
  wire n_2697_v;
  wire n_2706_v;
  wire n_634_v;
  wire n_2707_v;
  wire n_1011_v;
  wire n_2708_v;
  wire n_2741_v;
  wire n_1197_v;
  wire _t2_v;
  wire n_2326_v;
  wire n_1803_v;
  wire n_695_v;
  wire n_1236_v;
  wire m3_v;
  wire n_1348_v;
  wire n_1347_v;
  wire n_895_v;
  wire n_3484_v;
  wire n_1795_v;
  wire n_1798_v;
  wire n_1796_v;
  wire n_1799_v;
  wire n_890_v;
  wire n_3486_v;
  wire n_1797_v;
  wire n_1800_v;
  wire n_2333_v;
  wire n_3482_v;
  wire n_2336_v;
  wire n_3483_v;
  wire n_2332_v;
  wire n_3485_v;
  wire n_2334_v;
  wire n_2328_v;
  wire n_1787_v;
  wire n_782_v;
  wire n_3417_v;
  wire n_1495_v;
  wire n_484_v;
  wire n_780_v;
  wire n_3418_v;
  wire n_2725_v;
  wire n_2731_v;
  wire n_2726_v;
  wire n_2736_v;
  wire n_2727_v;
  wire n_2732_v;
  wire n_2728_v;
  wire n_2733_v;
  wire n_2729_v;
  wire n_2734_v;
  wire n_2730_v;
  wire n_2735_v;
  wire n_2017_v;
  wire n_793_v;
  wire n_82_v;
  wire n_1293_v;
  wire n_72_v;
  wire n_1402_v;
  wire n_406_v;
  wire n_2719_v;
  wire n_2742_v;
  wire n_1289_v;
  wire n_270_v;
  wire n_1108_v;
  wire n_1642_v;
  wire n_546_v;
  wire n_2043_v;
  wire n_1635_v;
  wire n_599_v;
  wire n_2709_v;
  wire n_2755_v;
  wire n_2710_v;
  wire n_2743_v;
  wire n_2711_v;
  wire n_2744_v;
  wire n_2712_v;
  wire n_2745_v;
  wire n_2713_v;
  wire n_2746_v;
  wire n_2714_v;
  wire n_2747_v;
  wire n_2749_v;
  wire n_2748_v;
  wire n_2342_v;
  wire n_3487_v;
  wire n_2750_v;
  wire n_2756_v;
  wire n_2716_v;
  wire n_2757_v;
  wire n_2717_v;
  wire n_2758_v;
  wire n_2752_v;
  wire n_2751_v;
  wire n_357_v;
  wire n_374_v;
  wire n_2753_v;
  wire n_2754_v;
  wire n_2718_v;
  wire n_2759_v;
  wire n_1497_v;
  wire n_330_v;
  wire n_46_v;
  wire ab5_v;
  wire ab6_v;
  wire ab7_v;
  wire ab8_v;
  wire ab9_v;
  wire ab10_v;
  wire ab11_v;
  wire ab12_v;
  wire ab13_v;
  wire ab14_v;
  wire ab15_v;
  wire n_1403_v;
  wire n_387_v;
  wire n_262_v;
  wire n_1426_v;
  wire n_1222_v;
  wire n_1229_v;
  wire n_233_v;
  wire n_135_v;
  wire n_1436_v;
  wire n_825_v;
  wire n_1433_v;
  wire n_1442_v;
  wire n_268_v;
  wire n_470_v;
  wire n_400_v;
  wire n_1435_v;
  wire n_826_v;
  wire n_1164_v;
  wire n_403_v;
  wire n_1456_v;
  wire n_424_v;
  wire n_1448_v;
  wire n_1465_v;
  wire n_191_v;
  wire n_1437_v;
  wire n_828_v;
  wire n_1210_v;
  wire n_361_v;
  wire n_1444_v;
  wire n_261_v;
  wire n_417_v;
  wire n_1463_v;
  wire n_413_v;
  wire n_459_v;
  wire n_1458_v;
  wire n_488_v;
  wire n_1445_v;
  wire n_1446_v;
  wire n_398_v;
  wire n_442_v;
  wire n_464_v;
  wire n_446_v;
  wire n_272_v;
  wire n_1467_v;
  wire n_349_v;
  wire n_273_v;
  wire n_1454_v;
  wire n_350_v;
  wire n_423_v;
  wire n_1459_v;
  wire n_427_v;
  wire n_468_v;
  wire n_391_v;
  wire n_432_v;
  wire n_457_v;
  wire n_1453_v;
  wire n_425_v;
  wire n_322_v;
  wire n_458_v;
  wire n_439_v;
  wire n_1450_v;
  wire n_449_v;
  wire n_409_v;
  wire n_1457_v;
  wire n_193_v;
  wire n_421_v;
  wire n_1461_v;
  wire n_428_v;
  wire n_1447_v;
  wire n_1091_v;
  wire n_469_v;
  wire n_422_v;
  wire n_401_v;
  wire n_453_v;
  wire n_1432_v;
  wire n_454_v;
  wire n_1438_v;
  wire n_1460_v;
  wire n_178_v;
  wire n_1246_v;
  wire n_1142_v;
  wire n_1425_v;
  wire n_1107_v;
  wire n_1100_v;
  wire n_1470_v;
  wire n_183_v;
  wire n_478_v;
  wire n_450_v;
  wire n_447_v;
  wire n_1233_v;
  wire n_184_v;
  wire n_1211_v;
  wire n_1215_v;
  wire n_1167_v;
  wire n_1474_v;
  wire n_1234_v;
  wire n_335_v;
  wire n_1057_v;
  wire n_249_v;
  wire n_236_v;
  wire n_1180_v;
  wire n_218_v;
  wire n_1102_v;
  wire n_76_v;
  wire n_1041_v;
  wire n_227_v;
  wire n_187_v;
  wire n_1237_v;
  wire n_200_v;
  wire n_1235_v;
  wire n_1147_v;
  wire n_1238_v;
  wire n_1213_v;
  wire n_53_v;
  wire n_289_v;
  wire n_104_v;
  wire n_1449_v;
  wire n_1089_v;
  wire n_202_v;
  wire n_1464_v;
  wire n_309_v;
  wire n_156_v;
  wire n_492_v;
  wire n_1476_v;
  wire n_1240_v;
  wire n_171_v;
  wire n_466_v;
  wire n_1477_v;
  wire n_1479_v;
  wire n_345_v;
  wire n_462_v;
  wire n_1469_v;
  wire n_463_v;
  wire n_467_v;
  wire n_441_v;
  wire n_1490_v;
  wire n_435_v;
  wire n_1489_v;
  wire n_430_v;
  wire n_1484_v;
  wire n_491_v;
  wire n_415_v;
  wire n_1486_v;
  wire n_1472_v;
  wire n_1468_v;
  wire n_1452_v;
  wire n_1493_v;
  wire n_1480_v;
  wire n_1475_v;
  wire n_1478_v;
  wire n_405_v;
  wire n_1494_v;
  wire n_1487_v;
  wire n_444_v;
  wire n_1483_v;
  wire n_404_v;
  wire n_1485_v;
  wire n_605_v;
  wire n_461_v;
  wire n_1481_v;
  wire n_1429_v;
  wire n_1488_v;
  wire n_455_v;
  wire n_1049_v;
  wire n_433_v;
  wire n_1255_v;
  wire n_352_v;
  wire n_1496_v;
  wire n_1244_v;
  wire n_186_v;
  wire n_1257_v;
  wire n_102_v;
  wire n_1109_v;
  wire n_1087_v;
  wire n_474_v;
  wire n_1491_v;
  wire n_1259_v;
  wire n_237_v;
  wire n_1250_v;
  wire n_1254_v;
  wire n_109_v;
  wire n_471_v;
  wire n_3014_v;
  wire n_174_v;
  wire n_245_v;
  wire n_231_v;
  wire n_1253_v;
  wire n_1262_v;
  wire n_1267_v;
  wire n_477_v;
  wire n_1501_v;
  wire n_476_v;
  wire n_182_v;
  wire n_74_v;
  wire n_1258_v;
  wire n_1499_v;
  wire n_1504_v;
  wire n_1083_v;
  wire n_1230_v;
  wire n_1273_v;
  wire n_1503_v;
  wire n_324_v;
  wire n_434_v;
  wire n_1500_v;
  wire n_1502_v;
  wire n_1260_v;
  wire n_229_v;
  wire n_1509_v;
  wire n_1274_v;
  wire n_1111_v;
  wire n_1508_v;
  wire n_487_v;
  wire n_271_v;
  wire n_323_v;
  wire n_1261_v;
  wire n_1266_v;
  wire n_1506_v;
  wire n_355_v;
  wire n_366_v;
  wire n_489_v;
  wire n_448_v;
  wire n_1231_v;
  wire n_296_v;
  wire n_1251_v;
  wire n_1263_v;
  wire n_1264_v;
  wire n_353_v;
  wire n_483_v;
  wire n_334_v;
  wire n_219_v;
  wire n_315_v;
  wire n_1512_v;
  wire n_1513_v;
  wire n_493_v;
  wire n_338_v;
  wire n_320_v;
  wire n_325_v;
  wire n_317_v;
  wire n_336_v;
  wire n_318_v;
  wire n_313_v;
  wire n_1516_v;
  wire n_52_v;
  wire n_290_v;
  wire n_363_v;
  wire n_495_v;
  wire n_198_v;
  wire n_497_v;
  wire n_473_v;
  wire n_1522_v;
  wire n_498_v;
  wire n_1521_v;
  wire n_1538_v;
  wire n_482_v;
  wire n_1519_v;
  wire n_501_v;
  wire n_1268_v;
  wire n_1272_v;
  wire n_63_v;
  wire n_1525_v;
  wire n_1539_v;
  wire n_1269_v;
  wire n_207_v;
  wire n_1114_v;
  wire n_112_v;
  wire n_300_v;
  wire n_206_v;
  wire n_1278_v;
  wire n_1084_v;
  wire n_1517_v;
  wire n_524_v;
  wire n_1256_v;
  wire n_201_v;
  wire n_514_v;
  wire n_1520_v;
  wire n_1540_v;
  wire n_365_v;
  wire n_287_v;
  wire n_1297_v;
  wire n_1524_v;
  wire n_504_v;
  wire n_205_v;
  wire n_1277_v;
  wire n_164_v;
  wire n_79_v;
  wire n_1116_v;
  wire n_1265_v;
  wire n_116_v;
  wire n_1545_v;
  wire n_460_v;
  wire n_1574_v;
  wire n_1527_v;
  wire n_1536_v;
  wire n_521_v;
  wire n_1543_v;
  wire n_1572_v;
  wire n_1549_v;
  wire n_1551_v;
  wire n_1534_v;
  wire n_1571_v;
  wire n_1537_v;
  wire n_542_v;
  wire n_213_v;
  wire n_1547_v;
  wire n_1594_v;
  wire n_1555_v;
  wire n_1591_v;
  wire n_1059_v;
  wire n_1055_v;
  wire n_1299_v;
  wire n_1279_v;
  wire n_1239_v;
  wire n_511_v;
  wire n_522_v;
  wire n_1291_v;
  wire n_1588_v;
  wire n_1189_v;
  wire n_543_v;
  wire n_1284_v;
  wire n_1559_v;
  wire n_1595_v;
  wire n_1562_v;
  wire n_1563_v;
  wire n_1535_v;
  wire n_1581_v;
  wire n_1564_v;
  wire n_1566_v;
  wire n_517_v;
  wire n_503_v;
  wire n_1548_v;
  wire n_1596_v;
  wire n_1528_v;
  wire n_1568_v;
  wire n_1587_v;
  wire n_91_v;
  wire n_1125_v;
  wire n_527_v;
  wire n_529_v;
  wire n_540_v;
  wire n_1567_v;
  wire n_1598_v;
  wire n_1542_v;
  wire n_536_v;
  wire n_1570_v;
  wire n_1606_v;
  wire n_1575_v;
  wire n_1592_v;
  wire n_530_v;
  wire n_203_v;
  wire n_55_v;
  wire n_224_v;
  wire n_215_v;
  wire n_515_v;
  wire n_1081_v;
  wire n_1082_v;
  wire n_1290_v;
  wire n_1066_v;
  wire n_1121_v;
  wire n_123_v;
  wire n_117_v;
  wire n_520_v;
  wire n_114_v;
  wire n_1110_v;
  wire n_239_v;
  wire n_1122_v;
  wire n_537_v;
  wire n_1569_v;
  wire n_1600_v;
  wire n_1046_v;
  wire n_1298_v;
  wire n_234_v;
  wire n_1123_v;
  wire n_1557_v;
  wire n_1576_v;
  wire n_130_v;
  wire n_195_v;
  wire n_1578_v;
  wire n_1580_v;
  wire n_1584_v;
  wire n_538_v;
  wire n_512_v;
  wire n_1560_v;
  wire n_535_v;
  wire n_1541_v;
  wire n_1597_v;
  wire n_1577_v;
  wire n_333_v;
  wire n_1124_v;
  wire n_1132_v;
  wire n_1602_v;
  wire n_1583_v;
  wire n_508_v;
  wire n_555_v;
  wire n_1601_v;
  wire n_539_v;
  wire n_1605_v;
  wire n_1553_v;
  wire n_1608_v;
  wire n_578_v;
  wire n_568_v;
  wire n_314_v;
  wire n_1558_v;
  wire n_1561_v;
  wire n_532_v;
  wire n_1603_v;
  wire n_533_v;
  wire n_332_v;
  wire n_513_v;
  wire n_507_v;
  wire n_1610_v;
  wire n_1565_v;
  wire n_1148_v;
  wire n_547_v;
  wire n_1589_v;
  wire n_1633_v;
  wire n_554_v;
  wire n_1515_v;
  wire n_1623_v;
  wire n_1604_v;
  wire n_583_v;
  wire n_1609_v;
  wire n_1624_v;
  wire n_306_v;
  wire n_1622_v;
  wire n_1523_v;
  wire n_1618_v;
  wire n_1612_v;
  wire n_1619_v;
  wire n_1532_v;
  wire n_1611_v;
  wire n_550_v;
  wire n_559_v;
  wire n_1645_v;
  wire n_1629_v;
  wire n_1550_v;
  wire n_1613_v;
  wire n_573_v;
  wire n_121_v;
  wire n_505_v;
  wire n_1643_v;
  wire n_1614_v;
  wire n_577_v;
  wire n_592_v;
  wire n_1616_v;
  wire n_1585_v;
  wire n_1641_v;
  wire n_518_v;
  wire n_581_v;
  wire n_593_v;
  wire n_1646_v;
  wire n_563_v;
  wire n_1636_v;
  wire n_1282_v;
  wire n_1621_v;
  wire n_1648_v;
  wire n_1137_v;
  wire n_211_v;
  wire n_1630_v;
  wire n_1632_v;
  wire n_561_v;
  wire n_1067_v;
  wire n_1128_v;
  wire n_569_v;
  wire n_1637_v;
  wire n_1639_v;
  wire n_1115_v;
  wire n_1112_v;
  wire n_1647_v;
  wire n_1105_v;
  wire n_1106_v;
  wire n_1152_v;
  wire n_1151_v;
  wire n_1133_v;
  wire n_1306_v;
  wire n_1307_v;
  wire n_1134_v;
  wire n_1135_v;
  wire n_1146_v;
  wire n_242_v;
  wire n_1308_v;
  wire n_1144_v;
  wire n_1138_v;
  wire n_125_v;
  wire n_567_v;
  wire n_1140_v;
  wire n_1319_v;
  wire n_1296_v;
  wire n_1310_v;
  wire n_285_v;
  wire n_230_v;
  wire n_1150_v;
  wire n_1662_v;
  wire n_1652_v;
  wire n_226_v;
  wire n_1136_v;
  wire n_1654_v;
  wire n_1127_v;
  wire n_113_v;
  wire n_310_v;
  wire n_1321_v;
  wire n_1324_v;
  wire n_1668_v;
  wire n_571_v;
  wire n_1659_v;
  wire n_1660_v;
  wire n_566_v;
  wire n_1141_v;
  wire n_579_v;
  wire n_580_v;
  wire n_1650_v;
  wire n_1664_v;
  wire n_601_v;
  wire n_1663_v;
  wire n_1657_v;
  wire n_572_v;
  wire n_1655_v;
  wire n_1640_v;
  wire n_591_v;
  wire n_685_v;
  wire n_1666_v;
  wire n_598_v;
  wire n_584_v;
  wire n_1615_v;
  wire n_1667_v;
  wire n_1656_v;
  wire n_264_v;
  wire n_238_v;
  wire n_160_v;
  wire n_1669_v;
  wire n_1323_v;
  wire n_1326_v;
  wire n_1670_v;
  wire n_610_v;
  wire n_1673_v;
  wire n_1672_v;
  wire n_1684_v;
  wire n_609_v;
  wire n_594_v;
  wire n_1677_v;
  wire n_619_v;
  wire n_499_v;
  wire n_1671_v;
  wire n_1676_v;
  wire n_1687_v;
  wire n_1688_v;
  wire n_1331_v;
  wire n_1248_v;
  wire n_1697_v;
  wire n_1143_v;
  wire n_611_v;
  wire n_1315_v;
  wire n_620_v;
  wire n_1682_v;
  wire n_1685_v;
  wire n_1675_v;
  wire n_1703_v;
  wire n_1681_v;
  wire n_1696_v;
  wire n_1314_v;
  wire n_269_v;
  wire n_1329_v;
  wire n_255_v;
  wire n_208_v;
  wire n_1305_v;
  wire n_582_v;
  wire n_1322_v;
  wire n_1695_v;
  wire n_252_v;
  wire n_628_v;
  wire n_632_v;
  wire n_1716_v;
  wire n_519_v;
  wire n_1287_v;
  wire n_1304_v;
  wire n_298_v;
  wire ex_dehl_combined_v;
  wire n_1713_v;
  wire n_1708_v;
  wire n_606_v;
  wire n_1711_v;
  wire n_630_v;
  wire n_1705_v;
  wire n_1712_v;
  wire n_1706_v;
  wire n_1714_v;
  wire n_1715_v;
  wire n_1704_v;
  wire n_1758_v;
  wire n_1333_v;
  wire n_311_v;
  wire n_1325_v;
  wire n_246_v;
  wire n_308_v;
  wire n_1294_v;
  wire n_1153_v;
  wire n_253_v;
  wire n_217_v;
  wire n_1710_v;
  wire n_312_v;
  wire n_1749_v;
  wire n_1750_v;
  wire n_1752_v;
  wire n_1693_v;
  wire n_712_v;
  wire n_1678_v;
  wire n_1755_v;
  wire n_1723_v;
  wire n_756_v;
  wire n_1700_v;
  wire n_624_v;
  wire n_1724_v;
  wire n_1683_v;
  wire n_623_v;
  wire n_637_v;
  wire n_1759_v;
  wire n_1727_v;
  wire n_1728_v;
  wire n_1334_v;
  wire n_1285_v;
  wire n_1730_v;
  wire n_1731_v;
  wire n_1720_v;
  wire n_649_v;
  wire n_1718_v;
  wire n_1764_v;
  wire n_638_v;
  wire n_648_v;
  wire n_636_v;
  wire n_1732_v;
  wire n_635_v;
  wire n_1721_v;
  wire n_1756_v;
  wire n_1763_v;
  wire n_1757_v;
  wire n_1726_v;
  wire n_1729_v;
  wire n_1157_v;
  wire n_221_v;
  wire n_1158_v;
  wire n_1155_v;
  wire n_1337_v;
  wire n_1734_v;
  wire n_141_v;
  wire n_1735_v;
  wire n_295_v;
  wire n_1073_v;
  wire n_1159_v;
  wire n_1733_v;
  wire n_1725_v;
  wire n_1160_v;
  wire n_256_v;
  wire n_60_v;
  wire n_640_v;
  wire n_1760_v;
  wire n_1145_v;
  wire n_1163_v;
  wire n_1768_v;
  wire n_1767_v;
  wire n_642_v;
  wire n_1765_v;
  wire n_639_v;
  wire n_1772_v;
  wire n_1771_v;
  wire n_1774_v;
  wire n_534_v;
  wire n_1722_v;
  wire n_1719_v;
  wire n_1165_v;
  wire n_1776_v;
  wire n_1777_v;
  wire n_1778_v;
  wire n_1781_v;
  wire n_1162_v;
  wire n_1172_v;
  wire n_644_v;
  wire n_1782_v;
  wire n_1794_v;
  wire n_1780_v;
  wire n_1793_v;
  wire n_1754_v;
  wire n_1775_v;
  wire n_1791_v;
  wire n_650_v;
  wire n_724_v;
  wire n_1182_v;
  wire n_1169_v;
  wire n_1423_v;
  wire n_683_v;
  wire n_686_v;
  wire n_1792_v;
  wire n_1738_v;
  wire n_1739_v;
  wire n_1740_v;
  wire n_1741_v;
  wire n_1742_v;
  wire n_1743_v;
  wire n_1744_v;
  wire n_1745_v;
  wire n_1746_v;
  wire n_1747_v;
  wire n_145_v;
  wire n_1806_v;
  wire n_1342_v;
  wire n_1187_v;
  wire n_1173_v;
  wire n_260_v;
  wire n_1175_v;
  wire n_1176_v;
  wire n_281_v;
  wire n_1343_v;
  wire n_257_v;
  wire n_1345_v;
  wire n_151_v;
  wire n_297_v;
  wire n_302_v;
  wire n_303_v;
  wire n_1805_v;
  wire n_258_v;
  wire n_304_v;
  wire n_305_v;
  wire n_277_v;
  wire n_278_v;
  wire n_279_v;
  wire n_282_v;
  wire n_283_v;
  wire n_284_v;
  wire n_286_v;
  wire n_1349_v;
  wire n_691_v;
  wire n_694_v;
  wire n_1807_v;
  wire n_698_v;
  wire n_329_v;
  wire n_1174_v;
  wire n_690_v;
  wire n_1809_v;
  wire n_1810_v;
  wire n_1813_v;
  wire n_699_v;
  wire n_1835_v;
  wire n_1832_v;
  wire n_1839_v;
  wire n_316_v;
  wire n_337_v;
  wire n_319_v;
  wire n_288_v;
  wire n_339_v;
  wire n_1808_v;
  wire n_340_v;
  wire n_341_v;
  wire n_291_v;
  wire n_1830_v;
  wire n_1829_v;
  wire n_342_v;
  wire n_1828_v;
  wire n_294_v;
  wire n_331_v;
  wire n_1831_v;
  wire n_1784_v;
  wire n_343_v;
  wire n_711_v;
  wire n_1862_v;
  wire n_1811_v;
  wire n_737_v;
  wire n_1857_v;
  wire n_1858_v;
  wire n_710_v;
  wire n_1856_v;
  wire n_344_v;
  wire n_1802_v;
  wire n_1812_v;
  wire n_1836_v;
  wire n_299_v;
  wire n_1855_v;
  wire n_301_v;
  wire n_346_v;
  wire n_266_v;
  wire n_347_v;
  wire n_348_v;
  wire n_1840_v;
  wire n_1863_v;
  wire n_307_v;
  wire n_276_v;
  wire n_1837_v;
  wire n_280_v;
  wire n_321_v;
  wire n_354_v;
  wire n_1351_v;
  wire n_1350_v;
  wire n_1353_v;
  wire n_1861_v;
  wire n_1166_v;
  wire n_1864_v;
  wire n_1865_v;
  wire n_1866_v;
  wire n_1867_v;
  wire n_1355_v;
  wire n_1352_v;
  wire n_356_v;
  wire n_274_v;
  wire n_351_v;
  wire n_275_v;
  wire n_1882_v;
  wire n_1886_v;
  wire n_765_v;
  wire n_730_v;
  wire n_1357_v;
  wire n_1860_v;
  wire n_717_v;
  wire n_736_v;
  wire n_364_v;
  wire n_727_v;
  wire n_1887_v;
  wire n_720_v;
  wire n_682_v;
  wire n_1908_v;
  wire n_764_v;
  wire n_729_v;
  wire n_768_v;
  wire n_292_v;
  wire n_1906_v;
  wire n_293_v;
  wire n_362_v;
  wire n_367_v;
  wire n_1930_v;
  wire n_1909_v;
  wire n_1904_v;
  wire n_368_v;
  wire n_1910_v;
  wire n_1907_v;
  wire n_1889_v;
  wire n_369_v;
  wire n_360_v;
  wire n_1356_v;
  wire n_402_v;
  wire n_372_v;
  wire n_1360_v;
  wire n_1789_v;
  wire n_1959_v;
  wire n_1943_v;
  wire n_1888_v;
  wire n_1944_v;
  wire n_1914_v;
  wire n_1937_v;
  wire n_1934_v;
  wire n_1931_v;
  wire n_758_v;
  wire n_1929_v;
  wire n_154_v;
  wire n_1938_v;
  wire n_1963_v;
  wire n_1960_v;
  wire n_748_v;
  wire n_1941_v;
  wire n_1967_v;
  wire n_1939_v;
  wire n_1188_v;
  wire n_1361_v;
  wire n_1363_v;
  wire n_751_v;
  wire n_1971_v;
  wire n_1972_v;
  wire n_1988_v;
  wire n_1859_v;
  wire n_1987_v;
  wire n_1992_v;
  wire n_773_v;
  wire n_377_v;
  wire n_358_v;
  wire n_1993_v;
  wire n_818_v;
  wire n_759_v;
  wire n_2011_v;
  wire n_1185_v;
  wire n_2012_v;
  wire n_1366_v;
  wire n_766_v;
  wire n_2013_v;
  wire n_2015_v;
  wire n_1995_v;
  wire n_1911_v;
  wire n_2016_v;
  wire n_1994_v;
  wire n_2018_v;
  wire n_2038_v;
  wire n_2035_v;
  wire n_778_v;
  wire n_2034_v;
  wire n_2033_v;
  wire n_97_v;
  wire n_2039_v;
  wire n_2060_v;
  wire n_2059_v;
  wire n_786_v;
  wire n_789_v;
  wire n_2090_v;
  wire n_2042_v;
  wire n_2065_v;
  wire n_2040_v;
  wire n_2067_v;
  wire n_2068_v;
  wire n_2085_v;
  wire n_251_v;
  wire n_2083_v;
  wire n_2088_v;
  wire n_2089_v;
  wire n_1367_v;
  wire n_1370_v;
  wire n_2113_v;
  wire n_2114_v;
  wire n_2093_v;
  wire n_2092_v;
  wire n_2118_v;
  wire n_2138_v;
  wire n_2135_v;
  wire n_152_v;
  wire n_2134_v;
  wire n_2133_v;
  wire n_2157_v;
  wire n_2156_v;
  wire n_811_v;
  wire n_842_v;
  wire n_2141_v;
  wire n_2159_v;
  wire n_2139_v;
  wire n_2161_v;
  wire n_2188_v;
  wire n_838_v;
  wire n_2162_v;
  wire n_2164_v;
  wire n_2165_v;
  wire n_2180_v;
  wire n_389_v;
  wire n_2187_v;
  wire n_854_v;
  wire n_2183_v;
  wire n_843_v;
  wire n_860_v;
  wire n_2213_v;
  wire n_2192_v;
  wire n_2193_v;
  wire n_2212_v;
  wire n_2220_v;
  wire n_2190_v;
  wire n_2216_v;
  wire n_2221_v;
  wire n_2222_v;
  wire n_1375_v;
  wire n_2195_v;
  wire n_865_v;
  wire n_855_v;
  wire n_2194_v;
  wire n_762_v;
  wire n_862_v;
  wire n_2218_v;
  wire n_2225_v;
  wire n_2228_v;
  wire n_866_v;
  wire n_872_v;
  wire n_2223_v;
  wire n_2252_v;
  wire n_2249_v;
  wire n_2219_v;
  wire n_2256_v;
  wire n_2255_v;
  wire n_2248_v;
  wire n_390_v;
  wire n_2246_v;
  wire n_882_v;
  wire n_876_v;
  wire n_2275_v;
  wire n_2274_v;
  wire n_869_v;
  wire n_1380_v;
  wire n_2276_v;
  wire n_2272_v;
  wire n_2277_v;
  wire n_2257_v;
  wire n_2278_v;
  wire n_2253_v;
  wire n_1190_v;
  wire n_2281_v;
  wire n_2282_v;
  wire n_2298_v;
  wire n_1048_v;
  wire n_1384_v;
  wire n_887_v;
  wire n_2297_v;
  wire n_2301_v;
  wire n_891_v;
  wire n_2303_v;
  wire n_2322_v;
  wire n_2331_v;
  wire n_905_v;
  wire n_2302_v;
  wire n_2323_v;
  wire n_2325_v;
  wire n_2324_v;
  wire n_153_v;
  wire n_1382_v;
  wire n_2329_v;
  wire n_2305_v;
  wire n_2327_v;
  wire n_894_v;
  wire n_2340_v;
  wire n_2304_v;
  wire n_2337_v;
  wire n_2335_v;
  wire n_2339_v;
  wire n_2341_v;
  wire n_2343_v;
  wire n_2365_v;
  wire n_2362_v;
  wire n_1389_v;
  wire n_1388_v;
  wire n_2361_v;
  wire n_2359_v;
  wire n_2370_v;
  wire n_912_v;
  wire n_904_v;
  wire n_2387_v;
  wire n_2385_v;
  wire n_1391_v;
  wire n_2358_v;
  wire n_394_v;
  wire n_2392_v;
  wire n_2368_v;
  wire n_2389_v;
  wire n_2394_v;
  wire n_2366_v;
  wire n_2369_v;
  wire n_2360_v;
  wire n_2400_v;
  wire n_2391_v;
  wire n_2399_v;
  wire n_2401_v;
  wire n_2402_v;
  wire n_2418_v;
  wire n_396_v;
  wire n_1395_v;
  wire n_1192_v;
  wire n_1396_v;
  wire n_1397_v;
  wire n_1179_v;
  wire n_2417_v;
  wire n_2422_v;
  wire n_1183_v;
  wire n_2425_v;
  wire n_932_v;
  wire n_919_v;
  wire n_2443_v;
  wire n_2423_v;
  wire n_2424_v;
  wire n_158_v;
  wire n_2446_v;
  wire n_1196_v;
  wire n_2447_v;
  wire n_1177_v;
  wire n_2448_v;
  wire n_167_v;
  wire n_2428_v;
  wire n_1200_v;
  wire n_1201_v;
  wire n_1195_v;
  wire n_2427_v;
  wire n_930_v;
  wire n_2449_v;
  wire n_2469_v;
  wire n_2466_v;
  wire n_1398_v;
  wire n_1054_v;
  wire n_381_v;
  wire n_1399_v;
  wire n_2465_v;
  wire n_2464_v;
  wire n_2474_v;
  wire n_2497_v;
  wire n_2475_v;
  wire n_1050_v;
  wire n_2495_v;
  wire n_2490_v;
  wire n_416_v;
  wire n_2472_v;
  wire n_2493_v;
  wire n_940_v;
  wire n_2503_v;
  wire n_2501_v;
  wire n_2502_v;
  wire n_2505_v;
  wire n_2473_v;
  wire n_2507_v;
  wire n_955_v;
  wire n_942_v;
  wire n_1052_v;
  wire n_2470_v;
  wire n_2508_v;
  wire n_2513_v;
  wire n_2529_v;
  wire n_2512_v;
  wire n_2530_v;
  wire n_410_v;
  wire n_2528_v;
  wire n_2534_v;
  wire n_960_v;
  wire n_952_v;
  wire n_2510_v;
  wire n_2536_v;
  wire n_2558_v;
  wire n_2535_v;
  wire n_2559_v;
  wire n_420_v;
  wire n_2562_v;
  wire n_2531_v;
  wire n_2538_v;
  wire n_1404_v;
  wire n_2511_v;
  wire n_2566_v;
  wire n_971_v;
  wire n_2557_v;
  wire n_2567_v;
  wire n_2537_v;
  wire n_2572_v;
  wire n_2592_v;
  wire n_2589_v;
  wire n_411_v;
  wire n_1212_v;
  wire n_1406_v;
  wire n_967_v;
  wire n_1407_v;
  wire n_2588_v;
  wire n_2587_v;
  wire n_2595_v;
  wire n_2570_v;
  wire n_1199_v;
  wire n_2612_v;
  wire n_2611_v;
  wire n_2596_v;
  wire n_2614_v;
  wire n_419_v;
  wire n_2593_v;
  wire n_2619_v;
  wire n_2618_v;
  wire n_1409_v;
  wire n_1410_v;
  wire n_2635_v;
  wire n_2661_v;
  wire n_2634_v;
  wire n_2638_v;
  wire n_2660_v;
  wire n_1096_v;
  wire n_407_v;
  wire n_414_v;
  wire n_2640_v;
  wire n_2657_v;
  wire n_986_v;
  wire n_2669_v;
  wire n_2670_v;
  wire n_2666_v;
  wire n_2667_v;
  wire n_2668_v;
  wire n_2671_v;
  wire n_2672_v;
  wire n_2674_v;
  wire n_1414_v;
  wire n_2642_v;
  wire n_1415_v;
  wire n_1099_v;
  wire n_2679_v;
  wire n_426_v;
  wire n_1002_v;
  wire n_997_v;
  wire n_2675_v;
  wire n_2681_v;
  wire n_2684_v;
  wire n_1000_v;
  wire n_2678_v;
  wire n_429_v;
  wire n_2689_v;
  wire n_2676_v;
  wire n_2691_v;
  wire n_2690_v;
  wire n_1412_v;
  wire n_1006_v;
  wire n_1026_v;
  wire n_2694_v;
  wire n_2692_v;
  wire n_1417_v;
  wire n_2698_v;
  wire n_1416_v;
  wire n_1419_v;
  wire n_1421_v;
  wire n_1424_v;
  wire n_1012_v;
  wire n_1013_v;
  wire n_1021_v;
  wire n_1022_v;
  wire n_1023_v;
  wire n_1024_v;
  wire n_1025_v;
  wire n_1015_v;
  wire n_1016_v;
  wire n_1019_v;
  wire n_179_v;
  wire n_47_v;
  wire n_2715_v;
  wire n_2720_v;
  wire n_2721_v;
  wire n_2722_v;
  wire n_2723_v;
  wire n_2724_v;
  wire n_1101_v;
  wire n_431_v;
  wire n_243_v;
  wire n_1198_v;
  wire n_2737_v;
  wire n_2738_v;
  wire n_2739_v;
  wire n_2740_v;
  wire n_1422_v;
  wire n_437_v;
  wire n_438_v;
  wire n_1420_v;
  wire n_1427_v;
  wire n_443_v;
  wire n_445_v;
  wire n_1431_v;
  wire n_180_v;
  wire n_1219_v;
  wire n_1227_v;
  wire n_1010_v;
  wire n_399_v;
  wire n_1413_v;
  wire n_516_v;
  wire n_1761_v;
  wire n_523_v;
  wire n_1554_v;
  wire n_1544_v;
  wire n_1531_v;
  wire n_1530_v;
  wire n_1518_v;
  wire n_1311_v;
  wire n_1208_v;
  wire n_1205_v;
  wire n_1699_v;
  wire n_1275_v;
  wire n_1276_v;
  wire n_645_v;
  wire n_212_v;
  wire n_1281_v;
  wire n_235_v;
  wire n_440_v;
  wire n_472_v;
  wire n_1283_v;
  wire n_531_v;
  wire n_1582_v;
  wire n_3358_v;
  wire n_1573_v;
  wire n_556_v;
  wire n_585_v;
  wire n_819_v;
  wire n_510_v;
  wire n_1131_v;
  wire n_1552_v;
  wire n_506_v;
  wire n_1085_v;
  wire n_189_v;
  wire n_490_v;
  wire n_1224_v;
  wire n_1206_v;
  wire n_688_v;
  wire n_1443_v;
  wire n_1628_v;
  wire n_565_v;
  wire n_1556_v;
  wire n_564_v;
  wire n_1252_v;
  wire n_1694_v;
  wire n_1411_v;
  wire n_1139_v;
  wire n_496_v;
  wire n_1526_v;
  wire n_500_v;
  wire n_1529_v;
  wire n_1686_v;
  wire n_1698_v;
  wire n_1690_v;
  wire n_1546_v;
  wire n_622_v;
  wire n_1689_v;
  wire n_1692_v;
  wire n_621_v;
  wire n_1691_v;
  wire n_1942_v;

  spice_pin_input pin_8659(_reset, _reset_v, _reset_port_1);
  spice_pin_input pin_8660(_wait, _wait_v, _wait_port_1);
  spice_pin_input pin_8661(_int, _int_v, _int_port_1);
  spice_pin_input pin_8662(_nmi, _nmi_v, _nmi_port_1);
  spice_pin_input pin_8663(_busrq, _busrq_v, _busrq_port_1);
  spice_pin_input pin_8672(clk, clk_v, clk_port_403);

  spice_pin_output pin_8635(ab0, a(ab0_v));
  spice_pin_output pin_8636(ab1, a(ab1_v));
  spice_pin_output pin_8637(ab2, a(ab2_v));
  spice_pin_output pin_8638(ab3, a(ab3_v));
  spice_pin_output pin_8639(ab4, a(ab4_v));
  spice_pin_output pin_8640(ab5, a(ab5_v));
  spice_pin_output pin_8641(ab6, a(ab6_v));
  spice_pin_output pin_8642(ab7, a(ab7_v));
  spice_pin_output pin_8643(ab8, a(ab8_v));
  spice_pin_output pin_8644(ab9, a(ab9_v));
  spice_pin_output pin_8645(ab10, a(ab10_v));
  spice_pin_output pin_8646(ab11, a(ab11_v));
  spice_pin_output pin_8647(ab12, a(ab12_v));
  spice_pin_output pin_8648(ab13, a(ab13_v));
  spice_pin_output pin_8649(ab14, a(ab14_v));
  spice_pin_output pin_8650(ab15, a(ab15_v));
  spice_pin_output pin_8664(_m1, a(_m1_v));
  spice_pin_output pin_8665(_rd, a(_rd_v));
  spice_pin_output pin_8666(_wr, a(_wr_v));
  spice_pin_output pin_8667(_mreq, a(_mreq_v));
  spice_pin_output pin_8668(_iorq, a(_iorq_v));
  spice_pin_output pin_8669(_rfsh, a(_rfsh_v));
  spice_pin_output pin_8670(_halt, a(_halt_v));
  spice_pin_output pin_8671(_busak, a(_busak_v));

  spice_pin_bidirectional pin_8651(db0_i, db0_o, db0_t, db0_v, db0_port_3);
  spice_pin_bidirectional pin_8652(db1_i, db1_o, db1_t, db1_v, db1_port_3);
  spice_pin_bidirectional pin_8653(db2_i, db2_o, db2_t, db2_v, db2_port_3);
  spice_pin_bidirectional pin_8654(db3_i, db3_o, db3_t, db3_v, db3_port_3);
  spice_pin_bidirectional pin_8655(db4_i, db4_o, db4_t, db4_v, db4_port_3);
  spice_pin_bidirectional pin_8656(db5_i, db5_o, db5_t, db5_v, db5_port_3);
  spice_pin_bidirectional pin_8657(db6_i, db6_o, db6_t, db6_v, db6_port_3);
  spice_pin_bidirectional pin_8658(db7_i, db7_o, db7_t, db7_v, db7_port_3);

  spice_transistor_nmos_vdd t2067(v(vcc_v), n_791_v, n_791_port_0);
  spice_transistor_nmos_vdd t2074(v(vcc_v), n_703_v, n_703_port_0);
  spice_transistor_nmos_vdd t2077(v(vcc_v), n_907_v, n_907_port_0);
  spice_transistor_nmos_vdd t2081(n_170_v, db0_v, db0_port_0);
  spice_transistor_nmos_vdd t2085(n_383_v, db7_v, db7_port_0);
  spice_transistor_nmos_vdd t2090(n_250_v, db1_v, db1_port_0);
  spice_transistor_nmos_vdd t2094(n_1507_v, n_380_v, n_380_port_0);
  spice_transistor_nmos_vdd t2095(n_1507_v, n_480_v, n_480_port_0);
  spice_transistor_nmos_vdd t2096(n_1507_v, n_485_v, n_485_port_0);
  spice_transistor_nmos_vdd t2097(n_1507_v, n_486_v, n_486_port_0);
  spice_transistor_nmos_vdd t2099(v(vcc_v), n_713_v, n_713_port_0);
  spice_transistor_nmos_vdd t2103(v(vcc_v), n_917_v, n_917_port_0);
  spice_transistor_nmos_vdd t2110(v(vcc_v), n_798_v, n_798_port_0);
  spice_transistor_nmos_vdd t2116(n_1507_v, n_370_v, n_370_port_0);
  spice_transistor_nmos_vdd t2120(n_1507_v, n_196_v, n_196_port_0);
  spice_transistor_nmos_vdd t2121(n_1507_v, n_412_v, n_412_port_0);
  spice_transistor_nmos_vdd t2122(n_1507_v, n_138_v, n_138_port_0);
  spice_transistor_nmos_vdd t2146(n_2108_v, n_790_v, n_790_port_0);
  spice_transistor_nmos_vdd t2148(v(vcc_v), n_922_v, n_922_port_0);
  spice_transistor_nmos_vdd t2159(v(vcc_v), n_806_v, n_806_port_0);
  spice_transistor_nmos_vdd t2176(n_2397_v, n_2338_v, n_2338_port_0);
  spice_transistor_nmos_vdd t2186(v(vcc_v), n_933_v, n_933_port_0);
  spice_transistor_nmos_vdd t2193(v(vcc_v), n_714_v, n_714_port_0);
  spice_transistor_nmos_vdd t2194(n_733_v, db6_v, db6_port_0);
  spice_transistor_nmos_vdd t2213(n_1379_v, n_248_v, n_248_port_0);
  spice_transistor_nmos_vdd t2228(n_1905_v, n_528_v, n_528_port_0);
  spice_transistor_nmos_vdd t2230(v(vcc_v), n_810_v, n_810_port_0);
  spice_transistor_nmos_vdd t2233(v(vcc_v), n_936_v, n_936_port_0);
  spice_transistor_nmos_vdd t2238(v(vcc_v), n_731_v, n_731_port_0);
  spice_transistor_nmos_vdd t2240(n_1707_v, n_616_v, n_616_port_0);
  spice_transistor_nmos_vdd t2246(n_821_v, n_944_v, n_944_port_0);
  spice_transistor_nmos_vdd t2251(n_2140_v, n_716_v, n_716_port_0);
  spice_transistor_nmos_vdd t2255(n_832_v, n_947_v, n_947_port_0);
  spice_transistor_nmos_vdd t2258(v(vcc_v), n_953_v, n_953_port_0);
  spice_transistor_nmos_vdd t2269(v(vcc_v), n_841_v, n_841_port_0);
  spice_transistor_nmos_vdd t2281(n_452_v, db2_v, db2_port_0);
  spice_transistor_nmos_vdd t2295(n_821_v, n_845_v, n_845_port_0);
  spice_transistor_nmos_vdd t2298(v(vcc_v), n_958_v, n_958_port_0);
  spice_transistor_nmos_vdd t2304(v(vcc_v), n_846_v, n_846_port_0);
  spice_transistor_nmos_vdd t2318(v(vcc_v), n_739_v, n_739_port_0);
  spice_transistor_nmos_vdd t2321(n_832_v, n_850_v, n_850_port_0);
  spice_transistor_nmos_vdd t2336(v(vcc_v), n_969_v, n_969_port_0);
  spice_transistor_nmos_vdd t2352(v(vcc_v), n_863_v, n_863_port_0);
  spice_transistor_nmos_vdd t2358(n_859_v, db5_v, db5_port_0);
  spice_transistor_nmos_vdd t2364(n_1940_v, n_526_v, n_526_port_0);
  spice_transistor_nmos_vdd t2374(n_978_v, db3_v, db3_port_0);
  spice_transistor_nmos_vdd t2380(v(vcc_v), n_749_v, n_749_port_0);
  spice_transistor_nmos_vdd t2398(v(vcc_v), n_974_v, n_974_port_0);
  spice_transistor_nmos_vdd t2402(n_2563_v, n_2504_v, n_2504_port_0);
  spice_transistor_nmos_vdd t2424(n_821_v, n_966_v, n_966_port_0);
  spice_transistor_nmos_vdd t2426(v(vcc_v), n_982_v, n_982_port_0);
  spice_transistor_nmos_vdd t2443(v(vcc_v), n_871_v, n_871_port_0);
  spice_transistor_nmos_vdd t2453(v(vcc_v), n_752_v, n_752_port_0);
  spice_transistor_nmos_vdd t2456(v(vcc_v), n_984_v, n_984_port_0);
  spice_transistor_nmos_vdd t2479(n_832_v, n_993_v, n_993_port_0);
  spice_transistor_nmos_vdd t2490(n_2247_v, n_2211_v, n_2211_port_0);
  spice_transistor_nmos_vdd t2492(v(vcc_v), n_884_v, n_884_port_0);
  spice_transistor_nmos_vdd t2493(v(vcc_v), n_998_v, n_998_port_0);
  spice_transistor_nmos_vdd t2517(v(vcc_v), n_774_v, n_774_port_0);
  spice_transistor_nmos_vdd t2532(v(vcc_v), n_885_v, n_885_port_0);
  spice_transistor_nmos_vdd t2559(n_2686_v, n_816_v, n_816_port_0);
  spice_transistor_nmos_vdd t2574(n_821_v, n_897_v, n_897_port_0);
  spice_transistor_nmos_vdd t2575(v(vcc_v), n_901_v, n_901_port_0);
  spice_transistor_nmos_vdd t2582(n_832_v, n_899_v, n_899_port_0);
  spice_transistor_nmos_vdd t2595(n_1787_v, n_697_v, n_697_port_0);
  spice_transistor_nmos_vdd t2597(v(vcc_v), n_777_v, n_777_port_0);
  spice_transistor_nmos_vdd t2683(n_1011_v, db4_v, db4_port_0);
  spice_transistor_nmos_gnd t2697(n_1439_v, db2_v, db2_port_1);
  spice_transistor_nmos_gnd t2719(n_1207_v, db0_v, db0_port_1);
  spice_transistor_nmos_gnd t2773(v(n_1232_v), n_190_v, n_190_port_0);
  spice_transistor_nmos_gnd t3395(v(n_1300_v), n_1302_v, n_1302_port_0);
  spice_transistor_nmos_gnd t3586(v(n_241_v), n_1332_v, n_1332_port_1);
  spice_transistor_nmos_gnd t3669(n_1685_v, n_616_v, n_616_port_1);
  spice_transistor_nmos_gnd t3780(n_1336_v, db1_v, db1_port_2);
  spice_transistor_nmos_gnd t3816(n_1753_v, db6_v, db6_port_1);
  spice_transistor_nmos_gnd t3903(n_637_v, n_647_v, n_647_port_0);
  spice_transistor_nmos_gnd t3936(v(n_58_v), n_1043_v, n_1043_port_1);
  spice_transistor_nmos_gnd t4101(n_637_v, n_701_v, n_701_port_0);
  spice_transistor_nmos_gnd t4102(n_1755_v, n_697_v, n_697_port_1);
  spice_transistor_nmos_gnd t4154(v(n_1814_v), reg_pcl0_v, reg_pcl0_port_0);
  spice_transistor_nmos_gnd t4155(v(n_1815_v), reg_r0_v, reg_r0_port_0);
  spice_transistor_nmos_gnd t4156(v(n_1816_v), reg_z0_v, reg_z0_port_0);
  spice_transistor_nmos_gnd t4157(v(n_1817_v), reg_spl0_v, reg_spl0_port_0);
  spice_transistor_nmos_gnd t4158(v(n_1818_v), reg_iyl0_v, reg_iyl0_port_0);
  spice_transistor_nmos_gnd t4159(v(n_1819_v), reg_ixl0_v, reg_ixl0_port_0);
  spice_transistor_nmos_gnd t4160(v(n_1820_v), reg_e0_v, reg_e0_port_0);
  spice_transistor_nmos_gnd t4161(v(n_1821_v), reg_ee0_v, reg_ee0_port_0);
  spice_transistor_nmos_gnd t4162(v(n_1822_v), reg_l0_v, reg_l0_port_0);
  spice_transistor_nmos_gnd t4163(v(n_1823_v), reg_ll0_v, reg_ll0_port_0);
  spice_transistor_nmos_gnd t4164(v(n_1824_v), reg_c0_v, reg_c0_port_0);
  spice_transistor_nmos_gnd t4165(v(n_1825_v), reg_cc0_v, reg_cc0_port_0);
  spice_transistor_nmos_gnd t4166(v(n_1826_v), reg_ff0_v, reg_ff0_port_0);
  spice_transistor_nmos_gnd t4167(v(n_1827_v), reg_f0_v, reg_f0_port_0);
  spice_transistor_nmos_gnd t4172(v(reg_pcl0_v), n_1814_v, n_1814_port_1);
  spice_transistor_nmos_gnd t4173(v(reg_r0_v), n_1815_v, n_1815_port_1);
  spice_transistor_nmos_gnd t4174(v(reg_z0_v), n_1816_v, n_1816_port_1);
  spice_transistor_nmos_gnd t4175(v(reg_spl0_v), n_1817_v, n_1817_port_1);
  spice_transistor_nmos_gnd t4176(v(reg_iyl0_v), n_1818_v, n_1818_port_1);
  spice_transistor_nmos_gnd t4177(v(reg_ixl0_v), n_1819_v, n_1819_port_1);
  spice_transistor_nmos_gnd t4178(v(reg_e0_v), n_1820_v, n_1820_port_1);
  spice_transistor_nmos_gnd t4179(v(reg_ee0_v), n_1821_v, n_1821_port_1);
  spice_transistor_nmos_gnd t4180(v(reg_l0_v), n_1822_v, n_1822_port_1);
  spice_transistor_nmos_gnd t4181(v(reg_ll0_v), n_1823_v, n_1823_port_1);
  spice_transistor_nmos_gnd t4182(v(reg_c0_v), n_1824_v, n_1824_port_1);
  spice_transistor_nmos_gnd t4183(v(reg_cc0_v), n_1825_v, n_1825_port_1);
  spice_transistor_nmos_gnd t4184(v(reg_ff0_v), n_1826_v, n_1826_port_1);
  spice_transistor_nmos_gnd t4185(v(reg_f0_v), n_1827_v, n_1827_port_1);
  spice_transistor_nmos_gnd t4240(n_1855_v, n_545_v, n_545_port_4);
  spice_transistor_nmos_gnd t4277(n_1882_v, n_528_v, n_528_port_1);
  spice_transistor_nmos_gnd t4290(v(reg_pcl1_v), n_1890_v, n_1890_port_0);
  spice_transistor_nmos_gnd t4291(v(reg_r1_v), n_1891_v, n_1891_port_0);
  spice_transistor_nmos_gnd t4293(v(reg_z1_v), n_1892_v, n_1892_port_0);
  spice_transistor_nmos_gnd t4294(v(reg_spl1_v), n_1893_v, n_1893_port_0);
  spice_transistor_nmos_gnd t4295(v(reg_iyl1_v), n_1894_v, n_1894_port_0);
  spice_transistor_nmos_gnd t4296(v(reg_ixl1_v), n_1895_v, n_1895_port_0);
  spice_transistor_nmos_gnd t4297(v(reg_e1_v), n_1896_v, n_1896_port_0);
  spice_transistor_nmos_gnd t4298(v(reg_ee1_v), n_1897_v, n_1897_port_0);
  spice_transistor_nmos_gnd t4299(v(reg_l1_v), n_1898_v, n_1898_port_0);
  spice_transistor_nmos_gnd t4300(v(reg_ll1_v), n_1899_v, n_1899_port_0);
  spice_transistor_nmos_gnd t4301(v(reg_c1_v), n_1900_v, n_1900_port_0);
  spice_transistor_nmos_gnd t4302(v(reg_cc1_v), n_1901_v, n_1901_port_0);
  spice_transistor_nmos_gnd t4303(v(reg_ff1_v), n_1902_v, n_1902_port_0);
  spice_transistor_nmos_gnd t4304(v(reg_f1_v), n_1903_v, n_1903_port_0);
  spice_transistor_nmos_gnd t4312(v(n_1890_v), reg_pcl1_v, reg_pcl1_port_1);
  spice_transistor_nmos_gnd t4313(v(n_1891_v), reg_r1_v, reg_r1_port_1);
  spice_transistor_nmos_gnd t4315(v(n_1892_v), reg_z1_v, reg_z1_port_1);
  spice_transistor_nmos_gnd t4316(v(n_1893_v), reg_spl1_v, reg_spl1_port_1);
  spice_transistor_nmos_gnd t4317(v(n_1894_v), reg_iyl1_v, reg_iyl1_port_1);
  spice_transistor_nmos_gnd t4318(v(n_1895_v), reg_ixl1_v, reg_ixl1_port_1);
  spice_transistor_nmos_gnd t4319(v(n_1896_v), reg_e1_v, reg_e1_port_1);
  spice_transistor_nmos_gnd t4320(v(n_1897_v), reg_ee1_v, reg_ee1_port_1);
  spice_transistor_nmos_gnd t4321(v(n_1898_v), reg_l1_v, reg_l1_port_1);
  spice_transistor_nmos_gnd t4322(v(n_1899_v), reg_ll1_v, reg_ll1_port_1);
  spice_transistor_nmos_gnd t4323(v(n_1900_v), reg_c1_v, reg_c1_port_1);
  spice_transistor_nmos_gnd t4324(v(n_1901_v), reg_cc1_v, reg_cc1_port_1);
  spice_transistor_nmos_gnd t4325(v(n_1902_v), reg_ff1_v, reg_ff1_port_1);
  spice_transistor_nmos_gnd t4326(v(n_1903_v), reg_f1_v, reg_f1_port_1);
  spice_transistor_nmos_gnd t4369(n_736_v, n_726_v, n_726_port_1);
  spice_transistor_nmos_gnd t4453(v(n_1915_v), reg_pcl2_v, reg_pcl2_port_0);
  spice_transistor_nmos_gnd t4454(v(n_1916_v), reg_r2_v, reg_r2_port_0);
  spice_transistor_nmos_gnd t4455(v(n_1917_v), reg_z2_v, reg_z2_port_0);
  spice_transistor_nmos_gnd t4456(v(n_1918_v), reg_spl2_v, reg_spl2_port_0);
  spice_transistor_nmos_gnd t4457(v(n_1919_v), reg_iyl2_v, reg_iyl2_port_0);
  spice_transistor_nmos_gnd t4458(v(n_1920_v), reg_ixl2_v, reg_ixl2_port_0);
  spice_transistor_nmos_gnd t4459(v(n_1921_v), reg_e2_v, reg_e2_port_0);
  spice_transistor_nmos_gnd t4460(v(n_1922_v), reg_ee2_v, reg_ee2_port_0);
  spice_transistor_nmos_gnd t4461(v(n_1923_v), reg_l2_v, reg_l2_port_0);
  spice_transistor_nmos_gnd t4462(v(n_1924_v), reg_ll2_v, reg_ll2_port_0);
  spice_transistor_nmos_gnd t4463(v(n_1925_v), reg_c2_v, reg_c2_port_0);
  spice_transistor_nmos_gnd t4464(v(n_1926_v), reg_cc2_v, reg_cc2_port_0);
  spice_transistor_nmos_gnd t4465(v(n_1927_v), reg_ff2_v, reg_ff2_port_0);
  spice_transistor_nmos_gnd t4466(v(n_1928_v), reg_f2_v, reg_f2_port_0);
  spice_transistor_nmos_gnd t4474(v(reg_pcl2_v), n_1915_v, n_1915_port_1);
  spice_transistor_nmos_gnd t4475(v(reg_r2_v), n_1916_v, n_1916_port_1);
  spice_transistor_nmos_gnd t4476(v(reg_z2_v), n_1917_v, n_1917_port_1);
  spice_transistor_nmos_gnd t4477(v(reg_spl2_v), n_1918_v, n_1918_port_1);
  spice_transistor_nmos_gnd t4478(v(reg_iyl2_v), n_1919_v, n_1919_port_1);
  spice_transistor_nmos_gnd t4479(v(reg_ixl2_v), n_1920_v, n_1920_port_1);
  spice_transistor_nmos_gnd t4480(v(reg_e2_v), n_1921_v, n_1921_port_1);
  spice_transistor_nmos_gnd t4481(v(reg_ee2_v), n_1922_v, n_1922_port_1);
  spice_transistor_nmos_gnd t4482(v(reg_l2_v), n_1923_v, n_1923_port_1);
  spice_transistor_nmos_gnd t4483(v(reg_ll2_v), n_1924_v, n_1924_port_1);
  spice_transistor_nmos_gnd t4484(v(reg_c2_v), n_1925_v, n_1925_port_1);
  spice_transistor_nmos_gnd t4485(v(reg_cc2_v), n_1926_v, n_1926_port_1);
  spice_transistor_nmos_gnd t4486(v(reg_ff2_v), n_1927_v, n_1927_port_1);
  spice_transistor_nmos_gnd t4487(v(reg_f2_v), n_1928_v, n_1928_port_1);
  spice_transistor_nmos_gnd t4528(n_1960_v, n_526_v, n_526_port_3);
  spice_transistor_nmos_gnd t4595(n_1987_v, n_770_v, n_770_port_2);
  spice_transistor_nmos_gnd t4607(v(reg_pcl3_v), n_1996_v, n_1996_port_0);
  spice_transistor_nmos_gnd t4608(v(reg_r3_v), n_1997_v, n_1997_port_0);
  spice_transistor_nmos_gnd t4610(v(reg_z3_v), n_1998_v, n_1998_port_0);
  spice_transistor_nmos_gnd t4611(v(reg_spl3_v), n_1999_v, n_1999_port_0);
  spice_transistor_nmos_gnd t4612(v(reg_iyl3_v), n_2000_v, n_2000_port_0);
  spice_transistor_nmos_gnd t4613(v(reg_ixl3_v), n_2001_v, n_2001_port_0);
  spice_transistor_nmos_gnd t4614(v(reg_e3_v), n_2002_v, n_2002_port_0);
  spice_transistor_nmos_gnd t4615(v(reg_ee3_v), n_2003_v, n_2003_port_0);
  spice_transistor_nmos_gnd t4616(v(reg_l3_v), n_2004_v, n_2004_port_0);
  spice_transistor_nmos_gnd t4617(v(reg_ll3_v), n_2005_v, n_2005_port_0);
  spice_transistor_nmos_gnd t4618(v(reg_c3_v), n_2006_v, n_2006_port_0);
  spice_transistor_nmos_gnd t4619(v(reg_cc3_v), n_2007_v, n_2007_port_0);
  spice_transistor_nmos_gnd t4620(v(reg_ff3_v), n_2008_v, n_2008_port_0);
  spice_transistor_nmos_gnd t4621(v(reg_f3_v), n_2009_v, n_2009_port_0);
  spice_transistor_nmos_gnd t4629(v(n_1996_v), reg_pcl3_v, reg_pcl3_port_1);
  spice_transistor_nmos_gnd t4630(v(n_1997_v), reg_r3_v, reg_r3_port_1);
  spice_transistor_nmos_gnd t4631(v(n_1998_v), reg_z3_v, reg_z3_port_1);
  spice_transistor_nmos_gnd t4632(v(n_1999_v), reg_spl3_v, reg_spl3_port_1);
  spice_transistor_nmos_gnd t4633(v(n_2000_v), reg_iyl3_v, reg_iyl3_port_1);
  spice_transistor_nmos_gnd t4634(v(n_2001_v), reg_ixl3_v, reg_ixl3_port_1);
  spice_transistor_nmos_gnd t4635(v(n_2002_v), reg_e3_v, reg_e3_port_1);
  spice_transistor_nmos_gnd t4636(v(n_2003_v), reg_ee3_v, reg_ee3_port_1);
  spice_transistor_nmos_gnd t4637(v(n_2004_v), reg_l3_v, reg_l3_port_1);
  spice_transistor_nmos_gnd t4638(v(n_2005_v), reg_ll3_v, reg_ll3_port_1);
  spice_transistor_nmos_gnd t4639(v(n_2006_v), reg_c3_v, reg_c3_port_1);
  spice_transistor_nmos_gnd t4640(v(n_2007_v), reg_cc3_v, reg_cc3_port_1);
  spice_transistor_nmos_gnd t4641(v(n_2008_v), reg_ff3_v, reg_ff3_port_1);
  spice_transistor_nmos_gnd t4642(v(n_2009_v), reg_f3_v, reg_f3_port_1);
  spice_transistor_nmos_gnd t4761(v(n_2019_v), reg_pcl4_v, reg_pcl4_port_0);
  spice_transistor_nmos_gnd t4762(v(n_2020_v), reg_r4_v, reg_r4_port_0);
  spice_transistor_nmos_gnd t4763(v(n_2021_v), reg_z4_v, reg_z4_port_0);
  spice_transistor_nmos_gnd t4764(v(n_2022_v), reg_spl4_v, reg_spl4_port_0);
  spice_transistor_nmos_gnd t4765(v(n_2023_v), reg_iyl4_v, reg_iyl4_port_0);
  spice_transistor_nmos_gnd t4766(v(n_2024_v), reg_ixl4_v, reg_ixl4_port_0);
  spice_transistor_nmos_gnd t4767(v(n_2025_v), reg_e4_v, reg_e4_port_0);
  spice_transistor_nmos_gnd t4768(v(n_2026_v), reg_ee4_v, reg_ee4_port_0);
  spice_transistor_nmos_gnd t4769(v(n_2027_v), reg_l4_v, reg_l4_port_0);
  spice_transistor_nmos_gnd t4770(v(n_2028_v), reg_ll4_v, reg_ll4_port_0);
  spice_transistor_nmos_gnd t4771(v(n_2029_v), reg_c4_v, reg_c4_port_0);
  spice_transistor_nmos_gnd t4772(v(n_2030_v), reg_cc4_v, reg_cc4_port_0);
  spice_transistor_nmos_gnd t4773(v(n_2031_v), reg_ff4_v, reg_ff4_port_0);
  spice_transistor_nmos_gnd t4774(v(n_2032_v), reg_f4_v, reg_f4_port_0);
  spice_transistor_nmos_gnd t4782(v(reg_pcl4_v), n_2019_v, n_2019_port_1);
  spice_transistor_nmos_gnd t4783(v(reg_r4_v), n_2020_v, n_2020_port_1);
  spice_transistor_nmos_gnd t4784(v(reg_z4_v), n_2021_v, n_2021_port_1);
  spice_transistor_nmos_gnd t4785(v(reg_spl4_v), n_2022_v, n_2022_port_1);
  spice_transistor_nmos_gnd t4786(v(reg_iyl4_v), n_2023_v, n_2023_port_1);
  spice_transistor_nmos_gnd t4787(v(reg_ixl4_v), n_2024_v, n_2024_port_1);
  spice_transistor_nmos_gnd t4788(v(reg_e4_v), n_2025_v, n_2025_port_1);
  spice_transistor_nmos_gnd t4789(v(reg_ee4_v), n_2026_v, n_2026_port_1);
  spice_transistor_nmos_gnd t4790(v(reg_l4_v), n_2027_v, n_2027_port_1);
  spice_transistor_nmos_gnd t4791(v(reg_ll4_v), n_2028_v, n_2028_port_1);
  spice_transistor_nmos_gnd t4792(v(reg_c4_v), n_2029_v, n_2029_port_1);
  spice_transistor_nmos_gnd t4793(v(reg_cc4_v), n_2030_v, n_2030_port_1);
  spice_transistor_nmos_gnd t4794(v(reg_ff4_v), n_2031_v, n_2031_port_1);
  spice_transistor_nmos_gnd t4795(v(reg_f4_v), n_2032_v, n_2032_port_1);
  spice_transistor_nmos_gnd t4831(n_2059_v, n_779_v, n_779_port_3);
  spice_transistor_nmos_gnd t4904(n_2083_v, n_790_v, n_790_port_1);
  spice_transistor_nmos_gnd t4916(v(reg_pcl5_v), n_2094_v, n_2094_port_0);
  spice_transistor_nmos_gnd t4917(v(reg_r5_v), n_2095_v, n_2095_port_0);
  spice_transistor_nmos_gnd t4919(v(reg_z5_v), n_2096_v, n_2096_port_0);
  spice_transistor_nmos_gnd t4920(v(reg_spl5_v), n_2097_v, n_2097_port_0);
  spice_transistor_nmos_gnd t4921(v(reg_iyl5_v), n_2098_v, n_2098_port_0);
  spice_transistor_nmos_gnd t4922(v(reg_ixl5_v), n_2099_v, n_2099_port_0);
  spice_transistor_nmos_gnd t4923(v(reg_e5_v), n_2100_v, n_2100_port_0);
  spice_transistor_nmos_gnd t4924(v(reg_ee5_v), n_2101_v, n_2101_port_0);
  spice_transistor_nmos_gnd t4925(v(reg_l5_v), n_2102_v, n_2102_port_0);
  spice_transistor_nmos_gnd t4926(v(reg_ll5_v), n_2103_v, n_2103_port_0);
  spice_transistor_nmos_gnd t4927(v(reg_c5_v), n_2104_v, n_2104_port_0);
  spice_transistor_nmos_gnd t4928(v(reg_cc5_v), n_2105_v, n_2105_port_0);
  spice_transistor_nmos_gnd t4929(v(reg_ff5_v), n_2106_v, n_2106_port_0);
  spice_transistor_nmos_gnd t4930(v(reg_f5_v), n_2107_v, n_2107_port_0);
  spice_transistor_nmos_gnd t4939(v(n_2094_v), reg_pcl5_v, reg_pcl5_port_1);
  spice_transistor_nmos_gnd t4940(v(n_2095_v), reg_r5_v, reg_r5_port_1);
  spice_transistor_nmos_gnd t4942(v(n_2096_v), reg_z5_v, reg_z5_port_1);
  spice_transistor_nmos_gnd t4943(v(n_2097_v), reg_spl5_v, reg_spl5_port_1);
  spice_transistor_nmos_gnd t4944(v(n_2098_v), reg_iyl5_v, reg_iyl5_port_1);
  spice_transistor_nmos_gnd t4945(v(n_2099_v), reg_ixl5_v, reg_ixl5_port_1);
  spice_transistor_nmos_gnd t4946(v(n_2100_v), reg_e5_v, reg_e5_port_1);
  spice_transistor_nmos_gnd t4947(v(n_2101_v), reg_ee5_v, reg_ee5_port_1);
  spice_transistor_nmos_gnd t4948(v(n_2102_v), reg_l5_v, reg_l5_port_1);
  spice_transistor_nmos_gnd t4949(v(n_2103_v), reg_ll5_v, reg_ll5_port_1);
  spice_transistor_nmos_gnd t4950(v(n_2104_v), reg_c5_v, reg_c5_port_1);
  spice_transistor_nmos_gnd t4951(v(n_2105_v), reg_cc5_v, reg_cc5_port_1);
  spice_transistor_nmos_gnd t4952(v(n_2106_v), reg_ff5_v, reg_ff5_port_1);
  spice_transistor_nmos_gnd t4953(v(n_2107_v), reg_f5_v, reg_f5_port_1);
  spice_transistor_nmos_gnd t5056(v(n_2119_v), reg_pcl6_v, reg_pcl6_port_0);
  spice_transistor_nmos_gnd t5057(v(n_2120_v), reg_r6_v, reg_r6_port_0);
  spice_transistor_nmos_gnd t5058(v(n_2121_v), reg_z6_v, reg_z6_port_0);
  spice_transistor_nmos_gnd t5059(v(n_2122_v), reg_spl6_v, reg_spl6_port_0);
  spice_transistor_nmos_gnd t5060(v(n_2123_v), reg_iyl6_v, reg_iyl6_port_0);
  spice_transistor_nmos_gnd t5061(v(n_2124_v), reg_ixl6_v, reg_ixl6_port_0);
  spice_transistor_nmos_gnd t5062(v(n_2125_v), reg_e6_v, reg_e6_port_0);
  spice_transistor_nmos_gnd t5063(v(n_2126_v), reg_ee6_v, reg_ee6_port_0);
  spice_transistor_nmos_gnd t5064(v(n_2127_v), reg_l6_v, reg_l6_port_0);
  spice_transistor_nmos_gnd t5065(v(n_2128_v), reg_ll6_v, reg_ll6_port_0);
  spice_transistor_nmos_gnd t5066(v(n_2129_v), reg_c6_v, reg_c6_port_0);
  spice_transistor_nmos_gnd t5067(v(n_2130_v), reg_cc6_v, reg_cc6_port_0);
  spice_transistor_nmos_gnd t5068(v(n_2131_v), reg_ff6_v, reg_ff6_port_0);
  spice_transistor_nmos_gnd t5069(v(n_2132_v), reg_f6_v, reg_f6_port_0);
  spice_transistor_nmos_gnd t5073(v(reg_pcl6_v), n_2119_v, n_2119_port_1);
  spice_transistor_nmos_gnd t5074(v(reg_r6_v), n_2120_v, n_2120_port_1);
  spice_transistor_nmos_gnd t5075(v(reg_z6_v), n_2121_v, n_2121_port_1);
  spice_transistor_nmos_gnd t5076(v(reg_spl6_v), n_2122_v, n_2122_port_1);
  spice_transistor_nmos_gnd t5077(v(reg_iyl6_v), n_2123_v, n_2123_port_1);
  spice_transistor_nmos_gnd t5078(v(reg_ixl6_v), n_2124_v, n_2124_port_1);
  spice_transistor_nmos_gnd t5079(v(reg_e6_v), n_2125_v, n_2125_port_1);
  spice_transistor_nmos_gnd t5080(v(reg_ee6_v), n_2126_v, n_2126_port_1);
  spice_transistor_nmos_gnd t5081(v(reg_l6_v), n_2127_v, n_2127_port_1);
  spice_transistor_nmos_gnd t5082(v(reg_ll6_v), n_2128_v, n_2128_port_1);
  spice_transistor_nmos_gnd t5083(v(reg_c6_v), n_2129_v, n_2129_port_1);
  spice_transistor_nmos_gnd t5084(v(reg_cc6_v), n_2130_v, n_2130_port_1);
  spice_transistor_nmos_gnd t5085(v(reg_ff6_v), n_2131_v, n_2131_port_1);
  spice_transistor_nmos_gnd t5086(v(reg_f6_v), n_2132_v, n_2132_port_1);
  spice_transistor_nmos_gnd t5103(n_2156_v, n_716_v, n_716_port_3);
  spice_transistor_nmos_gnd t5112(n_2158_v, db5_v, db5_port_1);
  spice_transistor_nmos_gnd t5145(n_2162_v, n_525_v, n_525_port_3);
  spice_transistor_nmos_gnd t5186(v(reg_pcl7_v), n_2196_v, n_2196_port_0);
  spice_transistor_nmos_gnd t5187(v(reg_r7_v), n_2197_v, n_2197_port_0);
  spice_transistor_nmos_gnd t5191(v(reg_z7_v), n_2198_v, n_2198_port_0);
  spice_transistor_nmos_gnd t5192(v(reg_spl7_v), n_2199_v, n_2199_port_0);
  spice_transistor_nmos_gnd t5193(v(reg_iyl7_v), n_2200_v, n_2200_port_0);
  spice_transistor_nmos_gnd t5194(v(reg_ixl7_v), n_2201_v, n_2201_port_0);
  spice_transistor_nmos_gnd t5195(v(reg_e7_v), n_2202_v, n_2202_port_0);
  spice_transistor_nmos_gnd t5196(v(reg_ee7_v), n_2203_v, n_2203_port_0);
  spice_transistor_nmos_gnd t5197(v(reg_l7_v), n_2204_v, n_2204_port_0);
  spice_transistor_nmos_gnd t5198(v(reg_ll7_v), n_2205_v, n_2205_port_0);
  spice_transistor_nmos_gnd t5199(v(reg_c7_v), n_2206_v, n_2206_port_0);
  spice_transistor_nmos_gnd t5200(v(reg_cc7_v), n_2207_v, n_2207_port_0);
  spice_transistor_nmos_gnd t5201(v(reg_ff7_v), n_2208_v, n_2208_port_0);
  spice_transistor_nmos_gnd t5202(v(reg_f7_v), n_2209_v, n_2209_port_0);
  spice_transistor_nmos_gnd t5215(v(n_2196_v), reg_pcl7_v, reg_pcl7_port_1);
  spice_transistor_nmos_gnd t5216(v(n_2197_v), reg_r7_v, reg_r7_port_1);
  spice_transistor_nmos_gnd t5219(v(n_2198_v), reg_z7_v, reg_z7_port_1);
  spice_transistor_nmos_gnd t5220(v(n_2199_v), reg_spl7_v, reg_spl7_port_1);
  spice_transistor_nmos_gnd t5221(v(n_2200_v), reg_iyl7_v, reg_iyl7_port_1);
  spice_transistor_nmos_gnd t5222(v(n_2201_v), reg_ixl7_v, reg_ixl7_port_1);
  spice_transistor_nmos_gnd t5223(v(n_2202_v), reg_e7_v, reg_e7_port_1);
  spice_transistor_nmos_gnd t5224(v(n_2203_v), reg_ee7_v, reg_ee7_port_1);
  spice_transistor_nmos_gnd t5225(v(n_2204_v), reg_l7_v, reg_l7_port_1);
  spice_transistor_nmos_gnd t5226(v(n_2205_v), reg_ll7_v, reg_ll7_port_1);
  spice_transistor_nmos_gnd t5227(v(n_2206_v), reg_c7_v, reg_c7_port_1);
  spice_transistor_nmos_gnd t5228(v(n_2207_v), reg_cc7_v, reg_cc7_port_1);
  spice_transistor_nmos_gnd t5229(v(n_2208_v), reg_ff7_v, reg_ff7_port_1);
  spice_transistor_nmos_gnd t5230(v(n_2209_v), reg_f7_v, reg_f7_port_1);
  spice_transistor_nmos_gnd t5289(n_1376_v, db7_v, db7_port_2);
  spice_transistor_nmos_gnd t5396(v(n_2232_v), reg_pch0_v, reg_pch0_port_0);
  spice_transistor_nmos_gnd t5397(v(n_2233_v), reg_i0_v, reg_i0_port_0);
  spice_transistor_nmos_gnd t5398(v(n_2234_v), reg_w0_v, reg_w0_port_0);
  spice_transistor_nmos_gnd t5399(v(n_2235_v), reg_sph0_v, reg_sph0_port_0);
  spice_transistor_nmos_gnd t5400(v(n_2236_v), reg_iyh0_v, reg_iyh0_port_0);
  spice_transistor_nmos_gnd t5401(v(n_2237_v), reg_ixh0_v, reg_ixh0_port_0);
  spice_transistor_nmos_gnd t5402(v(n_2238_v), reg_d0_v, reg_d0_port_0);
  spice_transistor_nmos_gnd t5403(v(n_2239_v), reg_dd0_v, reg_dd0_port_0);
  spice_transistor_nmos_gnd t5404(v(n_2240_v), reg_h0_v, reg_h0_port_0);
  spice_transistor_nmos_gnd t5405(v(n_2241_v), reg_hh0_v, reg_hh0_port_0);
  spice_transistor_nmos_gnd t5406(v(n_2242_v), reg_b0_v, reg_b0_port_0);
  spice_transistor_nmos_gnd t5407(v(n_2243_v), reg_bb0_v, reg_bb0_port_0);
  spice_transistor_nmos_gnd t5408(v(n_2244_v), reg_aa0_v, reg_aa0_port_0);
  spice_transistor_nmos_gnd t5409(v(n_2245_v), reg_a0_v, reg_a0_port_0);
  spice_transistor_nmos_gnd t5419(v(reg_pch0_v), n_2232_v, n_2232_port_1);
  spice_transistor_nmos_gnd t5420(v(reg_i0_v), n_2233_v, n_2233_port_1);
  spice_transistor_nmos_gnd t5421(v(reg_w0_v), n_2234_v, n_2234_port_1);
  spice_transistor_nmos_gnd t5422(v(reg_sph0_v), n_2235_v, n_2235_port_1);
  spice_transistor_nmos_gnd t5423(v(reg_iyh0_v), n_2236_v, n_2236_port_1);
  spice_transistor_nmos_gnd t5424(v(reg_ixh0_v), n_2237_v, n_2237_port_1);
  spice_transistor_nmos_gnd t5425(v(reg_d0_v), n_2238_v, n_2238_port_1);
  spice_transistor_nmos_gnd t5426(v(reg_dd0_v), n_2239_v, n_2239_port_1);
  spice_transistor_nmos_gnd t5427(v(reg_h0_v), n_2240_v, n_2240_port_1);
  spice_transistor_nmos_gnd t5428(v(reg_hh0_v), n_2241_v, n_2241_port_1);
  spice_transistor_nmos_gnd t5429(v(reg_b0_v), n_2242_v, n_2242_port_1);
  spice_transistor_nmos_gnd t5430(v(reg_bb0_v), n_2243_v, n_2243_port_1);
  spice_transistor_nmos_gnd t5431(v(reg_aa0_v), n_2244_v, n_2244_port_1);
  spice_transistor_nmos_gnd t5432(v(reg_a0_v), n_2245_v, n_2245_port_1);
  spice_transistor_nmos_gnd t5447(n_2219_v, n_2211_v, n_2211_port_3);
  spice_transistor_nmos_gnd t5452(n_388_v, n_248_v, n_248_port_25);
  spice_transistor_nmos_gnd t5534(v(reg_pch1_v), n_2306_v, n_2306_port_0);
  spice_transistor_nmos_gnd t5535(v(reg_i1_v), n_2307_v, n_2307_port_0);
  spice_transistor_nmos_gnd t5538(v(reg_w1_v), n_2308_v, n_2308_port_0);
  spice_transistor_nmos_gnd t5539(v(reg_sph1_v), n_2309_v, n_2309_port_0);
  spice_transistor_nmos_gnd t5540(v(reg_iyh1_v), n_2310_v, n_2310_port_0);
  spice_transistor_nmos_gnd t5541(v(reg_ixh1_v), n_2311_v, n_2311_port_0);
  spice_transistor_nmos_gnd t5542(v(reg_d1_v), n_2312_v, n_2312_port_0);
  spice_transistor_nmos_gnd t5543(v(reg_dd1_v), n_2313_v, n_2313_port_0);
  spice_transistor_nmos_gnd t5544(v(reg_h1_v), n_2314_v, n_2314_port_0);
  spice_transistor_nmos_gnd t5545(v(reg_hh1_v), n_2315_v, n_2315_port_0);
  spice_transistor_nmos_gnd t5546(v(reg_b1_v), n_2316_v, n_2316_port_0);
  spice_transistor_nmos_gnd t5547(v(reg_bb1_v), n_2317_v, n_2317_port_0);
  spice_transistor_nmos_gnd t5548(v(reg_aa1_v), n_2318_v, n_2318_port_0);
  spice_transistor_nmos_gnd t5549(v(reg_a1_v), n_2319_v, n_2319_port_0);
  spice_transistor_nmos_gnd t5556(v(n_2306_v), reg_pch1_v, reg_pch1_port_1);
  spice_transistor_nmos_gnd t5557(v(n_2307_v), reg_i1_v, reg_i1_port_1);
  spice_transistor_nmos_gnd t5558(v(n_2308_v), reg_w1_v, reg_w1_port_1);
  spice_transistor_nmos_gnd t5559(v(n_2309_v), reg_sph1_v, reg_sph1_port_1);
  spice_transistor_nmos_gnd t5560(v(n_2310_v), reg_iyh1_v, reg_iyh1_port_1);
  spice_transistor_nmos_gnd t5561(v(n_2311_v), reg_ixh1_v, reg_ixh1_port_1);
  spice_transistor_nmos_gnd t5562(v(n_2312_v), reg_d1_v, reg_d1_port_1);
  spice_transistor_nmos_gnd t5563(v(n_2313_v), reg_dd1_v, reg_dd1_port_1);
  spice_transistor_nmos_gnd t5564(v(n_2314_v), reg_h1_v, reg_h1_port_1);
  spice_transistor_nmos_gnd t5565(v(n_2315_v), reg_hh1_v, reg_hh1_port_1);
  spice_transistor_nmos_gnd t5566(v(n_2316_v), reg_b1_v, reg_b1_port_1);
  spice_transistor_nmos_gnd t5567(v(n_2317_v), reg_bb1_v, reg_bb1_port_1);
  spice_transistor_nmos_gnd t5568(v(n_2318_v), reg_aa1_v, reg_aa1_port_1);
  spice_transistor_nmos_gnd t5569(v(n_2319_v), reg_a1_v, reg_a1_port_1);
  spice_transistor_nmos_gnd t5698(v(n_2344_v), reg_pch2_v, reg_pch2_port_0);
  spice_transistor_nmos_gnd t5699(v(n_2345_v), reg_i2_v, reg_i2_port_0);
  spice_transistor_nmos_gnd t5700(v(n_2346_v), reg_w2_v, reg_w2_port_0);
  spice_transistor_nmos_gnd t5701(v(n_2347_v), reg_sph2_v, reg_sph2_port_0);
  spice_transistor_nmos_gnd t5702(v(n_2348_v), reg_iyh2_v, reg_iyh2_port_0);
  spice_transistor_nmos_gnd t5703(v(n_2349_v), reg_ixh2_v, reg_ixh2_port_0);
  spice_transistor_nmos_gnd t5704(v(n_2350_v), reg_d2_v, reg_d2_port_0);
  spice_transistor_nmos_gnd t5705(v(n_2351_v), reg_dd2_v, reg_dd2_port_0);
  spice_transistor_nmos_gnd t5706(v(n_2352_v), reg_h2_v, reg_h2_port_0);
  spice_transistor_nmos_gnd t5707(v(n_2353_v), reg_hh2_v, reg_hh2_port_0);
  spice_transistor_nmos_gnd t5708(v(n_2354_v), reg_b2_v, reg_b2_port_0);
  spice_transistor_nmos_gnd t5709(v(n_2355_v), reg_bb2_v, reg_bb2_port_0);
  spice_transistor_nmos_gnd t5710(v(n_2356_v), reg_aa2_v, reg_aa2_port_0);
  spice_transistor_nmos_gnd t5711(v(n_2357_v), reg_a2_v, reg_a2_port_0);
  spice_transistor_nmos_gnd t5724(v(reg_pch2_v), n_2344_v, n_2344_port_1);
  spice_transistor_nmos_gnd t5725(v(reg_i2_v), n_2345_v, n_2345_port_1);
  spice_transistor_nmos_gnd t5726(v(reg_w2_v), n_2346_v, n_2346_port_1);
  spice_transistor_nmos_gnd t5727(v(reg_sph2_v), n_2347_v, n_2347_port_1);
  spice_transistor_nmos_gnd t5728(v(reg_iyh2_v), n_2348_v, n_2348_port_1);
  spice_transistor_nmos_gnd t5729(v(reg_ixh2_v), n_2349_v, n_2349_port_1);
  spice_transistor_nmos_gnd t5730(v(reg_d2_v), n_2350_v, n_2350_port_1);
  spice_transistor_nmos_gnd t5731(v(reg_dd2_v), n_2351_v, n_2351_port_1);
  spice_transistor_nmos_gnd t5732(v(reg_h2_v), n_2352_v, n_2352_port_1);
  spice_transistor_nmos_gnd t5733(v(reg_hh2_v), n_2353_v, n_2353_port_1);
  spice_transistor_nmos_gnd t5734(v(reg_b2_v), n_2354_v, n_2354_port_1);
  spice_transistor_nmos_gnd t5735(v(reg_bb2_v), n_2355_v, n_2355_port_1);
  spice_transistor_nmos_gnd t5736(v(reg_aa2_v), n_2356_v, n_2356_port_1);
  spice_transistor_nmos_gnd t5737(v(reg_a2_v), n_2357_v, n_2357_port_1);
  spice_transistor_nmos_gnd t5874(v(reg_pch3_v), n_2429_v, n_2429_port_0);
  spice_transistor_nmos_gnd t5875(v(reg_i3_v), n_2430_v, n_2430_port_0);
  spice_transistor_nmos_gnd t5877(v(reg_w3_v), n_2431_v, n_2431_port_0);
  spice_transistor_nmos_gnd t5878(v(reg_sph3_v), n_2432_v, n_2432_port_0);
  spice_transistor_nmos_gnd t5879(v(reg_iyh3_v), n_2433_v, n_2433_port_0);
  spice_transistor_nmos_gnd t5880(v(reg_ixh3_v), n_2434_v, n_2434_port_0);
  spice_transistor_nmos_gnd t5881(v(reg_d3_v), n_2435_v, n_2435_port_0);
  spice_transistor_nmos_gnd t5882(v(reg_dd3_v), n_2436_v, n_2436_port_0);
  spice_transistor_nmos_gnd t5883(v(reg_h3_v), n_2437_v, n_2437_port_0);
  spice_transistor_nmos_gnd t5884(v(reg_hh3_v), n_2438_v, n_2438_port_0);
  spice_transistor_nmos_gnd t5885(v(reg_b3_v), n_2439_v, n_2439_port_0);
  spice_transistor_nmos_gnd t5886(v(reg_bb3_v), n_2440_v, n_2440_port_0);
  spice_transistor_nmos_gnd t5887(v(reg_aa3_v), n_2441_v, n_2441_port_0);
  spice_transistor_nmos_gnd t5888(v(reg_a3_v), n_2442_v, n_2442_port_0);
  spice_transistor_nmos_gnd t5897(n_2360_v, n_2338_v, n_2338_port_3);
  spice_transistor_nmos_gnd t5902(v(n_2429_v), reg_pch3_v, reg_pch3_port_1);
  spice_transistor_nmos_gnd t5903(v(n_2430_v), reg_i3_v, reg_i3_port_1);
  spice_transistor_nmos_gnd t5904(v(n_2431_v), reg_w3_v, reg_w3_port_1);
  spice_transistor_nmos_gnd t5905(v(n_2432_v), reg_sph3_v, reg_sph3_port_1);
  spice_transistor_nmos_gnd t5906(v(n_2433_v), reg_iyh3_v, reg_iyh3_port_1);
  spice_transistor_nmos_gnd t5907(v(n_2434_v), reg_ixh3_v, reg_ixh3_port_1);
  spice_transistor_nmos_gnd t5908(v(n_2435_v), reg_d3_v, reg_d3_port_1);
  spice_transistor_nmos_gnd t5909(v(n_2436_v), reg_dd3_v, reg_dd3_port_1);
  spice_transistor_nmos_gnd t5910(v(n_2437_v), reg_h3_v, reg_h3_port_1);
  spice_transistor_nmos_gnd t5911(v(n_2438_v), reg_hh3_v, reg_hh3_port_1);
  spice_transistor_nmos_gnd t5912(v(n_2439_v), reg_b3_v, reg_b3_port_1);
  spice_transistor_nmos_gnd t5913(v(n_2440_v), reg_bb3_v, reg_bb3_port_1);
  spice_transistor_nmos_gnd t5914(v(n_2441_v), reg_aa3_v, reg_aa3_port_1);
  spice_transistor_nmos_gnd t5915(v(n_2442_v), reg_a3_v, reg_a3_port_1);
  spice_transistor_nmos_gnd t6015(v(n_2450_v), reg_pch4_v, reg_pch4_port_0);
  spice_transistor_nmos_gnd t6016(v(n_2451_v), reg_i4_v, reg_i4_port_0);
  spice_transistor_nmos_gnd t6017(v(n_2452_v), reg_w4_v, reg_w4_port_0);
  spice_transistor_nmos_gnd t6018(v(n_2453_v), reg_sph4_v, reg_sph4_port_0);
  spice_transistor_nmos_gnd t6019(v(n_2454_v), reg_iyh4_v, reg_iyh4_port_0);
  spice_transistor_nmos_gnd t6020(v(n_2455_v), reg_ixh4_v, reg_ixh4_port_0);
  spice_transistor_nmos_gnd t6021(v(n_2456_v), reg_d4_v, reg_d4_port_0);
  spice_transistor_nmos_gnd t6022(v(n_2457_v), reg_dd4_v, reg_dd4_port_0);
  spice_transistor_nmos_gnd t6023(v(n_2458_v), reg_h4_v, reg_h4_port_0);
  spice_transistor_nmos_gnd t6024(v(n_2459_v), reg_hh4_v, reg_hh4_port_0);
  spice_transistor_nmos_gnd t6025(v(n_2460_v), reg_b4_v, reg_b4_port_0);
  spice_transistor_nmos_gnd t6026(v(n_2461_v), reg_bb4_v, reg_bb4_port_0);
  spice_transistor_nmos_gnd t6027(v(n_2462_v), reg_aa4_v, reg_aa4_port_0);
  spice_transistor_nmos_gnd t6028(v(n_2463_v), reg_a4_v, reg_a4_port_0);
  spice_transistor_nmos_gnd t6039(v(reg_pch4_v), n_2450_v, n_2450_port_1);
  spice_transistor_nmos_gnd t6040(v(reg_i4_v), n_2451_v, n_2451_port_1);
  spice_transistor_nmos_gnd t6041(v(reg_w4_v), n_2452_v, n_2452_port_1);
  spice_transistor_nmos_gnd t6042(v(reg_sph4_v), n_2453_v, n_2453_port_1);
  spice_transistor_nmos_gnd t6043(v(reg_iyh4_v), n_2454_v, n_2454_port_1);
  spice_transistor_nmos_gnd t6044(v(reg_ixh4_v), n_2455_v, n_2455_port_1);
  spice_transistor_nmos_gnd t6045(v(reg_d4_v), n_2456_v, n_2456_port_1);
  spice_transistor_nmos_gnd t6046(v(reg_dd4_v), n_2457_v, n_2457_port_1);
  spice_transistor_nmos_gnd t6047(v(reg_h4_v), n_2458_v, n_2458_port_1);
  spice_transistor_nmos_gnd t6048(v(reg_hh4_v), n_2459_v, n_2459_port_1);
  spice_transistor_nmos_gnd t6049(v(reg_b4_v), n_2460_v, n_2460_port_1);
  spice_transistor_nmos_gnd t6050(v(reg_bb4_v), n_2461_v, n_2461_port_1);
  spice_transistor_nmos_gnd t6051(v(reg_aa4_v), n_2462_v, n_2462_port_1);
  spice_transistor_nmos_gnd t6052(v(reg_a4_v), n_2463_v, n_2463_port_1);
  spice_transistor_nmos_gnd t6188(v(reg_pch5_v), n_2539_v, n_2539_port_0);
  spice_transistor_nmos_gnd t6189(v(reg_i5_v), n_2540_v, n_2540_port_0);
  spice_transistor_nmos_gnd t6192(v(reg_w5_v), n_2541_v, n_2541_port_0);
  spice_transistor_nmos_gnd t6193(v(reg_sph5_v), n_2542_v, n_2542_port_0);
  spice_transistor_nmos_gnd t6194(v(reg_iyh5_v), n_2543_v, n_2543_port_0);
  spice_transistor_nmos_gnd t6195(v(reg_ixh5_v), n_2544_v, n_2544_port_0);
  spice_transistor_nmos_gnd t6196(v(reg_d5_v), n_2545_v, n_2545_port_0);
  spice_transistor_nmos_gnd t6197(v(reg_dd5_v), n_2546_v, n_2546_port_0);
  spice_transistor_nmos_gnd t6198(v(reg_h5_v), n_2547_v, n_2547_port_0);
  spice_transistor_nmos_gnd t6199(v(reg_hh5_v), n_2548_v, n_2548_port_0);
  spice_transistor_nmos_gnd t6200(v(reg_b5_v), n_2549_v, n_2549_port_0);
  spice_transistor_nmos_gnd t6201(v(reg_bb5_v), n_2550_v, n_2550_port_0);
  spice_transistor_nmos_gnd t6202(v(reg_aa5_v), n_2551_v, n_2551_port_0);
  spice_transistor_nmos_gnd t6203(v(reg_a5_v), n_2552_v, n_2552_port_0);
  spice_transistor_nmos_gnd t6212(v(n_2539_v), reg_pch5_v, reg_pch5_port_1);
  spice_transistor_nmos_gnd t6213(v(n_2540_v), reg_i5_v, reg_i5_port_1);
  spice_transistor_nmos_gnd t6215(v(n_2541_v), reg_w5_v, reg_w5_port_1);
  spice_transistor_nmos_gnd t6216(v(n_2542_v), reg_sph5_v, reg_sph5_port_1);
  spice_transistor_nmos_gnd t6217(v(n_2543_v), reg_iyh5_v, reg_iyh5_port_1);
  spice_transistor_nmos_gnd t6218(v(n_2544_v), reg_ixh5_v, reg_ixh5_port_1);
  spice_transistor_nmos_gnd t6219(v(n_2545_v), reg_d5_v, reg_d5_port_1);
  spice_transistor_nmos_gnd t6220(v(n_2546_v), reg_dd5_v, reg_dd5_port_1);
  spice_transistor_nmos_gnd t6221(v(n_2547_v), reg_h5_v, reg_h5_port_1);
  spice_transistor_nmos_gnd t6222(v(n_2548_v), reg_hh5_v, reg_hh5_port_1);
  spice_transistor_nmos_gnd t6223(v(n_2549_v), reg_b5_v, reg_b5_port_1);
  spice_transistor_nmos_gnd t6224(v(n_2550_v), reg_bb5_v, reg_bb5_port_1);
  spice_transistor_nmos_gnd t6225(v(n_2551_v), reg_aa5_v, reg_aa5_port_1);
  spice_transistor_nmos_gnd t6226(v(n_2552_v), reg_a5_v, reg_a5_port_1);
  spice_transistor_nmos_gnd t6357(n_2511_v, n_2504_v, n_2504_port_3);
  spice_transistor_nmos_gnd t6380(v(n_2573_v), reg_pch6_v, reg_pch6_port_0);
  spice_transistor_nmos_gnd t6381(v(n_2574_v), reg_i6_v, reg_i6_port_0);
  spice_transistor_nmos_gnd t6382(v(n_2575_v), reg_w6_v, reg_w6_port_0);
  spice_transistor_nmos_gnd t6383(v(n_2576_v), reg_sph6_v, reg_sph6_port_0);
  spice_transistor_nmos_gnd t6384(v(n_2577_v), reg_iyh6_v, reg_iyh6_port_0);
  spice_transistor_nmos_gnd t6385(v(n_2578_v), reg_ixh6_v, reg_ixh6_port_0);
  spice_transistor_nmos_gnd t6386(v(n_2579_v), reg_d6_v, reg_d6_port_0);
  spice_transistor_nmos_gnd t6387(v(n_2580_v), reg_dd6_v, reg_dd6_port_0);
  spice_transistor_nmos_gnd t6388(v(n_2581_v), reg_h6_v, reg_h6_port_0);
  spice_transistor_nmos_gnd t6389(v(n_2582_v), reg_hh6_v, reg_hh6_port_0);
  spice_transistor_nmos_gnd t6390(v(n_2583_v), reg_b6_v, reg_b6_port_0);
  spice_transistor_nmos_gnd t6391(v(n_2584_v), reg_bb6_v, reg_bb6_port_0);
  spice_transistor_nmos_gnd t6392(v(n_2585_v), reg_aa6_v, reg_aa6_port_0);
  spice_transistor_nmos_gnd t6393(v(n_2586_v), reg_a6_v, reg_a6_port_0);
  spice_transistor_nmos_gnd t6399(v(reg_pch6_v), n_2573_v, n_2573_port_1);
  spice_transistor_nmos_gnd t6400(v(reg_i6_v), n_2574_v, n_2574_port_1);
  spice_transistor_nmos_gnd t6401(v(reg_w6_v), n_2575_v, n_2575_port_1);
  spice_transistor_nmos_gnd t6402(v(reg_sph6_v), n_2576_v, n_2576_port_1);
  spice_transistor_nmos_gnd t6403(v(reg_iyh6_v), n_2577_v, n_2577_port_1);
  spice_transistor_nmos_gnd t6404(v(reg_ixh6_v), n_2578_v, n_2578_port_1);
  spice_transistor_nmos_gnd t6405(v(reg_d6_v), n_2579_v, n_2579_port_1);
  spice_transistor_nmos_gnd t6406(v(reg_dd6_v), n_2580_v, n_2580_port_1);
  spice_transistor_nmos_gnd t6407(v(reg_h6_v), n_2581_v, n_2581_port_1);
  spice_transistor_nmos_gnd t6408(v(reg_hh6_v), n_2582_v, n_2582_port_1);
  spice_transistor_nmos_gnd t6409(v(reg_b6_v), n_2583_v, n_2583_port_1);
  spice_transistor_nmos_gnd t6410(v(reg_bb6_v), n_2584_v, n_2584_port_1);
  spice_transistor_nmos_gnd t6411(v(reg_aa6_v), n_2585_v, n_2585_port_1);
  spice_transistor_nmos_gnd t6412(v(reg_a6_v), n_2586_v, n_2586_port_1);
  spice_transistor_nmos_gnd t6468(n_2615_v, db3_v, db3_port_2);
  spice_transistor_nmos_gnd t6512(v(reg_pch7_v), n_2643_v, n_2643_port_0);
  spice_transistor_nmos_gnd t6513(v(reg_i7_v), n_2644_v, n_2644_port_0);
  spice_transistor_nmos_gnd t6515(v(reg_w7_v), n_2645_v, n_2645_port_0);
  spice_transistor_nmos_gnd t6516(v(reg_sph7_v), n_2646_v, n_2646_port_0);
  spice_transistor_nmos_gnd t6517(v(reg_iyh7_v), n_2647_v, n_2647_port_0);
  spice_transistor_nmos_gnd t6518(v(reg_ixh7_v), n_2648_v, n_2648_port_0);
  spice_transistor_nmos_gnd t6519(v(reg_d7_v), n_2649_v, n_2649_port_0);
  spice_transistor_nmos_gnd t6520(v(reg_dd7_v), n_2650_v, n_2650_port_0);
  spice_transistor_nmos_gnd t6521(v(reg_h7_v), n_2651_v, n_2651_port_0);
  spice_transistor_nmos_gnd t6522(v(reg_hh7_v), n_2652_v, n_2652_port_0);
  spice_transistor_nmos_gnd t6523(v(reg_b7_v), n_2653_v, n_2653_port_0);
  spice_transistor_nmos_gnd t6524(v(reg_bb7_v), n_2654_v, n_2654_port_0);
  spice_transistor_nmos_gnd t6525(v(reg_aa7_v), n_2655_v, n_2655_port_0);
  spice_transistor_nmos_gnd t6526(v(reg_a7_v), n_2656_v, n_2656_port_0);
  spice_transistor_nmos_gnd t6537(v(n_2643_v), reg_pch7_v, reg_pch7_port_1);
  spice_transistor_nmos_gnd t6538(v(n_2644_v), reg_i7_v, reg_i7_port_1);
  spice_transistor_nmos_gnd t6541(v(n_2645_v), reg_w7_v, reg_w7_port_1);
  spice_transistor_nmos_gnd t6542(v(n_2646_v), reg_sph7_v, reg_sph7_port_1);
  spice_transistor_nmos_gnd t6543(v(n_2647_v), reg_iyh7_v, reg_iyh7_port_1);
  spice_transistor_nmos_gnd t6544(v(n_2648_v), reg_ixh7_v, reg_ixh7_port_1);
  spice_transistor_nmos_gnd t6545(v(n_2649_v), reg_d7_v, reg_d7_port_1);
  spice_transistor_nmos_gnd t6546(v(n_2650_v), reg_dd7_v, reg_dd7_port_1);
  spice_transistor_nmos_gnd t6547(v(n_2651_v), reg_h7_v, reg_h7_port_1);
  spice_transistor_nmos_gnd t6548(v(n_2652_v), reg_hh7_v, reg_hh7_port_1);
  spice_transistor_nmos_gnd t6549(v(n_2653_v), reg_b7_v, reg_b7_port_1);
  spice_transistor_nmos_gnd t6550(v(n_2654_v), reg_bb7_v, reg_bb7_port_1);
  spice_transistor_nmos_gnd t6551(v(n_2655_v), reg_aa7_v, reg_aa7_port_1);
  spice_transistor_nmos_gnd t6552(v(n_2656_v), reg_a7_v, reg_a7_port_1);
  spice_transistor_nmos_gnd t6709(n_2676_v, n_816_v, n_816_port_4);
  spice_transistor_nmos_gnd t6781(n_2706_v, db4_v, db4_port_1);
  spice_transistor_nmos t7017(n_662_v, n_753_v, reg_e3_v, n_753_port_1, reg_e3_port_2);
  spice_transistor_nmos t7020(n_665_v, reg_ee3_v, n_753_v, reg_ee3_port_2, n_753_port_2);
  spice_transistor_nmos t7022(n_666_v, n_753_v, reg_l3_v, n_753_port_3, reg_l3_port_2);
  spice_transistor_nmos t7023(n_793_v, n_889_v, n_772_v, n_889_port_1, n_772_port_5);
  spice_transistor_nmos t7028(n_669_v, reg_ll3_v, n_753_v, reg_ll3_port_2, n_753_port_4);
  spice_transistor_nmos t7029(n_1799_v, n_901_v, n_2306_v, n_901_port_2, n_2306_port_2);
  spice_transistor_nmos t7030(n_1800_v, n_2307_v, n_901_v, n_2307_port_2, n_901_port_3);
  spice_transistor_nmos t7031(n_670_v, n_753_v, reg_c3_v, n_753_port_5, reg_c3_port_2);
  spice_transistor_nmos t7032(n_654_v, n_902_v, n_2308_v, n_902_port_0, n_2308_port_2);
  spice_transistor_nmos t7033(n_657_v, n_2309_v, n_902_v, n_2309_port_2, n_902_port_1);
  spice_transistor_nmos t7034(n_658_v, n_902_v, n_2310_v, n_902_port_2, n_2310_port_2);
  spice_transistor_nmos t7035(n_661_v, n_2311_v, n_902_v, n_2311_port_2, n_902_port_3);
  spice_transistor_nmos t7036(n_662_v, n_902_v, n_2312_v, n_902_port_4, n_2312_port_2);
  spice_transistor_nmos t7037(n_665_v, n_2313_v, n_902_v, n_2313_port_2, n_902_port_5);
  spice_transistor_nmos t7038(n_666_v, n_902_v, n_2314_v, n_902_port_6, n_2314_port_2);
  spice_transistor_nmos t7039(n_669_v, n_2315_v, n_902_v, n_2315_port_2, n_902_port_7);
  spice_transistor_nmos t7040(n_670_v, n_902_v, n_2316_v, n_902_port_8, n_2316_port_2);
  spice_transistor_nmos t7041(n_673_v, n_2317_v, n_902_v, n_2317_port_2, n_902_port_9);
  spice_transistor_nmos t7042(n_674_v, n_902_v, n_2318_v, n_902_port_10, n_2318_port_2);
  spice_transistor_nmos t7043(n_677_v, n_2319_v, n_902_v, n_2319_port_2, n_902_port_11);
  spice_transistor_nmos t7046(n_673_v, reg_cc3_v, n_753_v, reg_cc3_port_2, n_753_port_6);
  spice_transistor_nmos t7047(n_674_v, n_753_v, reg_ff3_v, n_753_port_7, reg_ff3_port_2);
  spice_transistor_nmos t7050(n_677_v, reg_f3_v, n_753_v, reg_f3_port_2, n_753_port_8);
  wire [`W-1:0] temp_12444;
  spice_transistor_nmos t7071(n_1994_v, a(n_1988_v), n_763_v, temp_12444, n_763_port_2);
  spice_transistor_nmos t7086(n_1799_v, n_907_v, n_2344_v, n_907_port_3, n_2344_port_2);
  spice_transistor_nmos t7087(n_1800_v, n_2345_v, n_907_v, n_2345_port_2, n_907_port_4);
  spice_transistor_nmos t7088(n_654_v, n_906_v, n_2346_v, n_906_port_0, n_2346_port_2);
  spice_transistor_nmos t7089(n_657_v, n_2347_v, n_906_v, n_2347_port_2, n_906_port_1);
  spice_transistor_nmos t7090(n_658_v, n_906_v, n_2348_v, n_906_port_2, n_2348_port_2);
  spice_transistor_nmos t7091(n_661_v, n_2349_v, n_906_v, n_2349_port_2, n_906_port_3);
  spice_transistor_nmos t7092(n_662_v, n_906_v, n_2350_v, n_906_port_4, n_2350_port_2);
  spice_transistor_nmos t7093(n_665_v, n_2351_v, n_906_v, n_2351_port_2, n_906_port_5);
  spice_transistor_nmos t7094(n_666_v, n_906_v, n_2352_v, n_906_port_6, n_2352_port_2);
  spice_transistor_nmos t7095(n_669_v, n_2353_v, n_906_v, n_2353_port_2, n_906_port_7);
  spice_transistor_nmos t7096(n_670_v, n_906_v, n_2354_v, n_906_port_8, n_2354_port_2);
  spice_transistor_nmos t7097(n_673_v, n_2355_v, n_906_v, n_2355_port_2, n_906_port_9);
  spice_transistor_nmos t7098(n_674_v, n_906_v, n_2356_v, n_906_port_10, n_2356_port_2);
  spice_transistor_nmos t7099(n_677_v, n_2357_v, n_906_v, n_2357_port_2, n_906_port_11);
  spice_transistor_nmos t7101(n_1785_v, n_907_v, n_906_v, n_907_port_5, n_906_port_13);
  wire [`W-1:0] temp_12445;
  spice_transistor_nmos t7110(n_2358_v, a(n_2340_v), n_908_v, temp_12445, n_908_port_1);
  wire [`W-1:0] temp_12446;
  spice_transistor_nmos t7111(n_1995_v, a(n_1971_v), n_769_v, temp_12446, n_769_port_1);
  spice_transistor_nmos t7133(n_735_v, n_783_v, n_889_v, n_783_port_5, n_889_port_2);
  spice_transistor_nmos t7137(n_750_v, n_772_v, n_528_v, n_772_port_6, n_528_port_3);
  wire [`W-1:0] temp_12447;
  spice_transistor_nmos t7142(n_2366_v, a(n_2362_v), n_913_v, temp_12447, n_913_port_0);
  wire [`W-1:0] temp_12448;
  spice_transistor_nmos t7147(n_1971_v, a(n_1995_v), n_769_v, temp_12448, n_769_port_2);
  wire [`W-1:0] temp_12449;
  spice_transistor_nmos t7149(n_1988_v, n_763_v, a(n_1994_v), n_763_port_3, temp_12449);
  wire [`W-1:0] temp_12450;
  spice_transistor_nmos t7151(n_2368_v, a(n_2365_v), n_915_v, temp_12450, n_915_port_2);
  spice_transistor_nmos t7156(n_1785_v, n_774_v, n_775_v, n_774_port_3, n_775_port_1);
  wire [`W-1:0] temp_12451;
  spice_transistor_nmos t7157(n_766_v, n_754_v, a(n_2011_v), n_754_port_1, temp_12451);
  wire [`W-1:0] temp_12452;
  spice_transistor_nmos t7168(n_2011_v, a(n_766_v), n_754_v, temp_12452, n_754_port_2);
  spice_transistor_nmos t7178(v(n_1061_v), n_2775_v, n_2776_v, n_2775_port_0, n_2776_port_0);
  spice_transistor_nmos t7179(n_643_v, n_889_v, n_755_v, n_889_port_3, n_755_port_5);
  wire [`W-1:0] temp_12453;
  spice_transistor_nmos t7181(n_2340_v, n_908_v, a(n_2358_v), n_908_port_2, temp_12453);
  spice_transistor_nmos t7197(n_1799_v, n_774_v, n_1996_v, n_774_port_4, n_1996_port_2);
  spice_transistor_nmos t7198(n_1800_v, n_1997_v, n_774_v, n_1997_port_2, n_774_port_5);
  spice_transistor_nmos t7199(n_654_v, n_775_v, n_1998_v, n_775_port_3, n_1998_port_2);
  spice_transistor_nmos t7200(n_657_v, n_1999_v, n_775_v, n_1999_port_2, n_775_port_4);
  spice_transistor_nmos t7201(n_658_v, n_775_v, n_2000_v, n_775_port_5, n_2000_port_2);
  spice_transistor_nmos t7202(n_661_v, n_2001_v, n_775_v, n_2001_port_2, n_775_port_6);
  spice_transistor_nmos t7203(n_662_v, n_775_v, n_2002_v, n_775_port_7, n_2002_port_2);
  spice_transistor_nmos t7204(n_665_v, n_2003_v, n_775_v, n_2003_port_2, n_775_port_8);
  spice_transistor_nmos t7205(n_666_v, n_775_v, n_2004_v, n_775_port_9, n_2004_port_2);
  spice_transistor_nmos t7206(n_669_v, n_2005_v, n_775_v, n_2005_port_2, n_775_port_10);
  spice_transistor_nmos t7207(n_670_v, n_775_v, n_2006_v, n_775_port_11, n_2006_port_2);
  spice_transistor_nmos t7208(n_673_v, n_2007_v, n_775_v, n_2007_port_2, n_775_port_12);
  wire [`W-1:0] temp_12454;
  spice_transistor_nmos t7209(n_2365_v, a(n_2368_v), n_915_v, temp_12454, n_915_port_3);
  spice_transistor_nmos t7210(n_674_v, n_775_v, n_2008_v, n_775_port_13, n_2008_port_2);
  spice_transistor_nmos t7212(n_677_v, n_2009_v, n_775_v, n_2009_port_2, n_775_port_14);
  spice_transistor_nmos t7219(n_1785_v, n_917_v, n_914_v, n_917_port_1, n_914_port_1);
  wire [`W-1:0] temp_12455;
  spice_transistor_nmos t7228(n_2362_v, n_913_v, a(n_2366_v), n_913_port_1, temp_12455);
  wire [`W-1:0] temp_12456;
  spice_transistor_nmos t7231(n_183_v, n_181_v, a(n_1239_v), n_181_port_4, temp_12456);
  wire [`W-1:0] temp_12457;
  spice_transistor_nmos t7240(n_636_v, n_647_v, a(n_1784_v), n_647_port_3, temp_12457);
  spice_transistor_nmos t7244(n_546_v, n_770_v, n_480_v, n_770_port_4, n_480_port_7);
  spice_transistor_nmos t7248(n_1799_v, n_917_v, reg_pch2_v, n_917_port_3, reg_pch2_port_2);
  spice_transistor_nmos t7249(n_1800_v, reg_i2_v, n_917_v, reg_i2_port_2, n_917_port_4);
  spice_transistor_nmos t7250(n_654_v, n_914_v, reg_w2_v, n_914_port_4, reg_w2_port_2);
  spice_transistor_nmos t7251(n_657_v, reg_sph2_v, n_914_v, reg_sph2_port_2, n_914_port_5);
  spice_transistor_nmos t7252(n_658_v, n_914_v, reg_iyh2_v, n_914_port_6, reg_iyh2_port_2);
  spice_transistor_nmos t7253(n_661_v, reg_ixh2_v, n_914_v, reg_ixh2_port_2, n_914_port_7);
  spice_transistor_nmos t7254(n_662_v, n_914_v, reg_d2_v, n_914_port_8, reg_d2_port_2);
  spice_transistor_nmos t7255(n_665_v, reg_dd2_v, n_914_v, reg_dd2_port_2, n_914_port_9);
  spice_transistor_nmos t7256(n_666_v, n_914_v, reg_h2_v, n_914_port_10, reg_h2_port_2);
  spice_transistor_nmos t7257(n_669_v, reg_hh2_v, n_914_v, reg_hh2_port_2, n_914_port_11);
  spice_transistor_nmos t7258(n_670_v, n_914_v, reg_b2_v, n_914_port_12, reg_b2_port_2);
  spice_transistor_nmos t7259(n_673_v, reg_bb2_v, n_914_v, reg_bb2_port_2, n_914_port_13);
  spice_transistor_nmos t7260(n_674_v, n_914_v, reg_aa2_v, n_914_port_14, reg_aa2_port_2);
  spice_transistor_nmos t7261(n_677_v, reg_a2_v, n_914_v, reg_a2_port_2, n_914_port_15);
  spice_transistor_nmos t7268(n_643_v, n_803_v, n_903_v, n_803_port_5, n_903_port_2);
  spice_transistor_nmos t7269(n_750_v, n_526_v, n_783_v, n_526_port_6, n_783_port_6);
  spice_transistor_nmos t7272(n_575_v, n_647_v, n_526_v, n_647_port_4, n_526_port_7);
  spice_transistor_nmos t7274(n_1799_v, n_777_v, n_2019_v, n_777_port_3, n_2019_port_2);
  spice_transistor_nmos t7275(n_1800_v, n_2020_v, n_777_v, n_2020_port_2, n_777_port_4);
  spice_transistor_nmos t7276(n_654_v, n_776_v, n_2021_v, n_776_port_0, n_2021_port_2);
  spice_transistor_nmos t7277(n_657_v, n_2022_v, n_776_v, n_2022_port_2, n_776_port_1);
  spice_transistor_nmos t7278(n_658_v, n_776_v, n_2023_v, n_776_port_2, n_2023_port_2);
  spice_transistor_nmos t7279(n_661_v, n_2024_v, n_776_v, n_2024_port_2, n_776_port_3);
  spice_transistor_nmos t7280(n_662_v, n_776_v, n_2025_v, n_776_port_4, n_2025_port_2);
  spice_transistor_nmos t7281(n_665_v, n_2026_v, n_776_v, n_2026_port_2, n_776_port_5);
  spice_transistor_nmos t7282(n_666_v, n_776_v, n_2027_v, n_776_port_6, n_2027_port_2);
  spice_transistor_nmos t7283(n_669_v, n_2028_v, n_776_v, n_2028_port_2, n_776_port_7);
  spice_transistor_nmos t7284(n_670_v, n_776_v, n_2029_v, n_776_port_8, n_2029_port_2);
  spice_transistor_nmos t7285(n_673_v, n_2030_v, n_776_v, n_2030_port_2, n_776_port_9);
  spice_transistor_nmos t7286(n_674_v, n_776_v, n_2031_v, n_776_port_10, n_2031_port_2);
  spice_transistor_nmos t7287(n_677_v, n_2032_v, n_776_v, n_2032_port_2, n_776_port_11);
  spice_transistor_nmos t7289(n_1785_v, n_777_v, n_776_v, n_777_port_5, n_776_port_13);
  spice_transistor_nmos t7311(n_735_v, n_903_v, n_836_v, n_903_port_3, n_836_port_5);
  spice_transistor_nmos t7322(n_1785_v, n_922_v, n_923_v, n_922_port_2, n_923_port_1);
  spice_transistor_nmos t7328(n_1799_v, n_922_v, reg_pch3_v, n_922_port_3, reg_pch3_port_2);
  spice_transistor_nmos t7331(n_1800_v, reg_i3_v, n_922_v, reg_i3_port_2, n_922_port_4);
  spice_transistor_nmos t7337(n_654_v, n_923_v, reg_w3_v, n_923_port_4, reg_w3_port_2);
  spice_transistor_nmos t7340(n_657_v, reg_sph3_v, n_923_v, reg_sph3_port_2, n_923_port_5);
  spice_transistor_nmos t7341(n_658_v, n_923_v, reg_iyh3_v, n_923_port_6, reg_iyh3_port_2);
  spice_transistor_nmos t7344(n_661_v, reg_ixh3_v, n_923_v, reg_ixh3_port_2, n_923_port_7);
  spice_transistor_nmos t7345(n_662_v, n_923_v, reg_d3_v, n_923_port_8, reg_d3_port_2);
  wire [`W-1:0] temp_12458;
  spice_transistor_nmos t7346(n_2040_v, a(n_2035_v), n_784_v, temp_12458, n_784_port_0);
  spice_transistor_nmos t7348(n_665_v, reg_dd3_v, n_923_v, reg_dd3_port_2, n_923_port_9);
  spice_transistor_nmos t7349(n_666_v, n_923_v, reg_h3_v, n_923_port_10, reg_h3_port_2);
  spice_transistor_nmos t7350(n_546_v, n_779_v, n_485_v, n_779_port_4, n_485_port_7);
  spice_transistor_nmos t7352(n_669_v, reg_hh3_v, n_923_v, reg_hh3_port_2, n_923_port_11);
  spice_transistor_nmos t7353(n_670_v, n_923_v, reg_b3_v, n_923_port_12, reg_b3_port_2);
  spice_transistor_nmos t7356(n_673_v, reg_bb3_v, n_923_v, reg_bb3_port_2, n_923_port_13);
  spice_transistor_nmos t7357(n_674_v, n_923_v, reg_aa3_v, n_923_port_14, reg_aa3_port_2);
  spice_transistor_nmos t7360(n_677_v, reg_a3_v, n_923_v, reg_a3_port_2, n_923_port_15);
  wire [`W-1:0] temp_12459;
  spice_transistor_nmos t7365(n_2042_v, a(n_2038_v), n_787_v, temp_12459, n_787_port_3);
  spice_transistor_nmos t7372(n_207_v, n_181_v, n_248_v, n_181_port_5, n_248_port_26);
  wire [`W-1:0] temp_12460;
  spice_transistor_nmos t7386(v(clk_v), a(n_1792_v), n_647_v, temp_12460, n_647_port_5);
  wire [`W-1:0] temp_12461;
  spice_transistor_nmos t7387(n_2427_v, a(n_2418_v), n_928_v, temp_12461, n_928_port_1);
  spice_transistor_nmos t7389(n_750_v, n_770_v, n_796_v, n_770_port_5, n_796_port_5);
  wire [`W-1:0] temp_12462;
  spice_transistor_nmos t7407(n_2428_v, a(n_2401_v), n_929_v, temp_12462, n_929_port_1);
  wire [`W-1:0] temp_12463;
  spice_transistor_nmos t7423(n_2038_v, a(n_2042_v), n_787_v, temp_12463, n_787_port_4);
  spice_transistor_nmos t7431(n_1785_v, n_791_v, n_785_v, n_791_port_1, n_785_port_1);
  spice_transistor_nmos t7433(n_546_v, n_790_v, n_486_v, n_790_port_3, n_486_port_6);
  wire [`W-1:0] temp_12464;
  spice_transistor_nmos t7439(n_2035_v, n_784_v, a(n_2040_v), n_784_port_1, temp_12464);
  spice_transistor_nmos t7447(n_793_v, n_808_v, n_903_v, n_808_port_5, n_903_port_5);
  wire [`W-1:0] temp_12465;
  spice_transistor_nmos t7450(n_2401_v, a(n_2428_v), n_929_v, temp_12465, n_929_port_2);
  wire [`W-1:0] temp_12466;
  spice_transistor_nmos t7452(n_2418_v, n_928_v, a(n_2427_v), n_928_port_2, temp_12466);
  spice_transistor_nmos t7459(n_1785_v, n_933_v, n_934_v, n_933_port_3, n_934_port_1);
  wire [`W-1:0] temp_12467;
  spice_transistor_nmos t7461(v(clk_v), a(n_2399_v), n_918_v, temp_12467, n_918_port_1);
  spice_transistor_nmos t7470(n_1799_v, n_791_v, reg_pcl4_v, n_791_port_3, reg_pcl4_port_2);
  spice_transistor_nmos t7471(n_1800_v, reg_r4_v, n_791_v, reg_r4_port_2, n_791_port_4);
  spice_transistor_nmos t7472(n_654_v, n_785_v, reg_z4_v, n_785_port_4, reg_z4_port_2);
  wire [`W-1:0] temp_12468;
  spice_transistor_nmos t7475(n_740_v, a(n_2423_v), n_918_v, temp_12468, n_918_port_3);
  spice_transistor_nmos t7476(n_657_v, reg_spl4_v, n_785_v, reg_spl4_port_2, n_785_port_5);
  spice_transistor_nmos t7477(n_658_v, n_785_v, reg_iyl4_v, n_785_port_6, reg_iyl4_port_2);
  spice_transistor_nmos t7478(n_820_v, n_918_v, n_903_v, n_918_port_4, n_903_port_8);
  spice_transistor_nmos t7480(n_661_v, reg_ixl4_v, n_785_v, reg_ixl4_port_2, n_785_port_7);
  spice_transistor_nmos t7481(n_662_v, n_785_v, reg_e4_v, n_785_port_8, reg_e4_port_2);
  spice_transistor_nmos t7482(n_665_v, reg_ee4_v, n_785_v, reg_ee4_port_2, n_785_port_9);
  spice_transistor_nmos t7483(n_666_v, n_785_v, reg_l4_v, n_785_port_10, reg_l4_port_2);
  spice_transistor_nmos t7484(n_646_v, n_2338_v, n_903_v, n_2338_port_5, n_903_port_10);
  spice_transistor_nmos t7485(n_669_v, reg_ll4_v, n_785_v, reg_ll4_port_2, n_785_port_11);
  spice_transistor_nmos t7486(n_670_v, n_785_v, reg_c4_v, n_785_port_12, reg_c4_port_2);
  spice_transistor_nmos t7487(n_673_v, reg_cc4_v, n_785_v, reg_cc4_port_2, n_785_port_13);
  spice_transistor_nmos t7489(n_674_v, n_785_v, reg_ff4_v, n_785_port_14, reg_ff4_port_2);
  spice_transistor_nmos t7490(n_677_v, reg_f4_v, n_785_v, reg_f4_port_2, n_785_port_15);
  spice_transistor_nmos t7495(n_1799_v, n_933_v, n_2429_v, n_933_port_4, n_2429_port_2);
  spice_transistor_nmos t7496(n_1800_v, n_2430_v, n_933_v, n_2430_port_2, n_933_port_5);
  spice_transistor_nmos t7497(n_654_v, n_934_v, n_2431_v, n_934_port_3, n_2431_port_2);
  spice_transistor_nmos t7498(n_657_v, n_2432_v, n_934_v, n_2432_port_2, n_934_port_4);
  spice_transistor_nmos t7499(n_658_v, n_934_v, n_2433_v, n_934_port_5, n_2433_port_2);
  spice_transistor_nmos t7500(n_661_v, n_2434_v, n_934_v, n_2434_port_2, n_934_port_6);
  spice_transistor_nmos t7501(n_662_v, n_934_v, n_2435_v, n_934_port_7, n_2435_port_2);
  spice_transistor_nmos t7502(n_665_v, n_2436_v, n_934_v, n_2436_port_2, n_934_port_8);
  spice_transistor_nmos t7503(n_666_v, n_934_v, n_2437_v, n_934_port_9, n_2437_port_2);
  spice_transistor_nmos t7504(n_669_v, n_2438_v, n_934_v, n_2438_port_2, n_934_port_10);
  spice_transistor_nmos t7505(n_670_v, n_934_v, n_2439_v, n_934_port_11, n_2439_port_2);
  spice_transistor_nmos t7506(n_673_v, n_2440_v, n_934_v, n_2440_port_2, n_934_port_12);
  spice_transistor_nmos t7507(n_674_v, n_934_v, n_2441_v, n_934_port_13, n_2441_port_2);
  spice_transistor_nmos t7508(n_677_v, n_2442_v, n_934_v, n_2442_port_2, n_934_port_14);
  spice_transistor_nmos t7530(n_1799_v, n_936_v, n_2450_v, n_936_port_3, n_2450_port_2);
  spice_transistor_nmos t7531(n_1800_v, n_2451_v, n_936_v, n_2451_port_2, n_936_port_4);
  spice_transistor_nmos t7532(n_654_v, n_935_v, n_2452_v, n_935_port_0, n_2452_port_2);
  spice_transistor_nmos t7533(n_657_v, n_2453_v, n_935_v, n_2453_port_2, n_935_port_1);
  spice_transistor_nmos t7534(n_658_v, n_935_v, n_2454_v, n_935_port_2, n_2454_port_2);
  spice_transistor_nmos t7535(n_661_v, n_2455_v, n_935_v, n_2455_port_2, n_935_port_3);
  spice_transistor_nmos t7536(n_662_v, n_935_v, n_2456_v, n_935_port_4, n_2456_port_2);
  spice_transistor_nmos t7537(n_665_v, n_2457_v, n_935_v, n_2457_port_2, n_935_port_5);
  spice_transistor_nmos t7538(n_666_v, n_935_v, n_2458_v, n_935_port_6, n_2458_port_2);
  spice_transistor_nmos t7539(n_669_v, n_2459_v, n_935_v, n_2459_port_2, n_935_port_7);
  spice_transistor_nmos t7540(n_670_v, n_935_v, n_2460_v, n_935_port_8, n_2460_port_2);
  spice_transistor_nmos t7541(n_673_v, n_2461_v, n_935_v, n_2461_port_2, n_935_port_9);
  spice_transistor_nmos t7542(n_674_v, n_935_v, n_2462_v, n_935_port_10, n_2462_port_2);
  spice_transistor_nmos t7543(n_677_v, n_2463_v, n_935_v, n_2463_port_2, n_935_port_11);
  spice_transistor_nmos t7545(n_1785_v, n_936_v, n_935_v, n_936_port_5, n_935_port_13);
  spice_transistor_nmos t7554(n_750_v, n_779_v, n_803_v, n_779_port_5, n_803_port_6);
  spice_transistor_nmos t7557(n_546_v, n_716_v, n_380_v, n_716_port_4, n_380_port_2);
  spice_transistor_nmos t7574(n_1785_v, n_798_v, n_799_v, n_798_port_2, n_799_port_1);
  wire [`W-1:0] temp_12469;
  spice_transistor_nmos t7579(n_2470_v, a(n_2466_v), n_948_v, temp_12469, n_948_port_0);
  spice_transistor_nmos t7582(n_1799_v, n_798_v, reg_pcl5_v, n_798_port_3, reg_pcl5_port_2);
  wire [`W-1:0] temp_12470;
  spice_transistor_nmos t7585(n_2473_v, a(n_2469_v), n_950_v, temp_12470, n_950_port_3);
  spice_transistor_nmos t7586(n_1800_v, reg_r5_v, n_798_v, reg_r5_port_2, n_798_port_4);
  spice_transistor_nmos t7591(n_654_v, n_799_v, reg_z5_v, n_799_port_4, reg_z5_port_2);
  spice_transistor_nmos t7594(n_657_v, reg_spl5_v, n_799_v, reg_spl5_port_2, n_799_port_5);
  spice_transistor_nmos t7595(n_658_v, n_799_v, reg_iyl5_v, n_799_port_6, reg_iyl5_port_2);
  spice_transistor_nmos t7598(n_661_v, reg_ixl5_v, n_799_v, reg_ixl5_port_2, n_799_port_7);
  spice_transistor_nmos t7599(n_662_v, n_799_v, reg_e5_v, n_799_port_8, reg_e5_port_2);
  spice_transistor_nmos t7602(n_665_v, reg_ee5_v, n_799_v, reg_ee5_port_2, n_799_port_9);
  spice_transistor_nmos t7603(n_666_v, n_799_v, reg_l5_v, n_799_port_10, reg_l5_port_2);
  wire [`W-1:0] temp_12471;
  spice_transistor_nmos t7606(n_740_v, n_944_v, a(n_940_v), n_944_port_2, temp_12471);
  wire [`W-1:0] temp_12472;
  spice_transistor_nmos t7608(n_740_v, a(n_2497_v), n_947_v, temp_12472, n_947_port_2);
  spice_transistor_nmos t7609(n_669_v, reg_ll5_v, n_799_v, reg_ll5_port_2, n_799_port_11);
  spice_transistor_nmos t7610(n_670_v, n_799_v, reg_c5_v, n_799_port_12, reg_c5_port_2);
  spice_transistor_nmos t7612(n_820_v, n_937_v, n_944_v, n_937_port_4, n_944_port_3);
  spice_transistor_nmos t7613(n_604_v, n_937_v, n_947_v, n_937_port_5, n_947_port_3);
  spice_transistor_nmos t7615(n_673_v, reg_cc5_v, n_799_v, reg_cc5_port_2, n_799_port_13);
  spice_transistor_nmos t7616(n_674_v, n_799_v, reg_ff5_v, n_799_port_14, reg_ff5_port_2);
  spice_transistor_nmos t7619(n_677_v, reg_f5_v, n_799_v, reg_f5_port_2, n_799_port_15);
  wire [`W-1:0] temp_12473;
  spice_transistor_nmos t7635(v(clk_v), n_947_v, a(n_2501_v), n_947_port_4, temp_12473);
  wire [`W-1:0] temp_12474;
  spice_transistor_nmos t7638(v(clk_v), n_944_v, a(n_2502_v), n_944_port_4, temp_12474);
  wire [`W-1:0] temp_12475;
  spice_transistor_nmos t7648(n_2092_v, a(n_2085_v), n_802_v, temp_12475, n_802_port_2);
  wire [`W-1:0] temp_12476;
  spice_transistor_nmos t7652(n_2469_v, a(n_2473_v), n_950_v, temp_12476, n_950_port_4);
  wire [`W-1:0] temp_12477;
  spice_transistor_nmos t7658(n_1758_v, a(n_635_v), n_697_v, temp_12477, n_697_port_3);
  spice_transistor_nmos t7662(n_1785_v, n_953_v, n_949_v, n_953_port_1, n_949_port_1);
  wire [`W-1:0] temp_12478;
  spice_transistor_nmos t7665(n_2466_v, n_948_v, a(n_2470_v), n_948_port_1, temp_12478);
  spice_transistor_nmos t7668(n_793_v, n_937_v, n_783_v, n_937_port_7, n_783_port_7);
  spice_transistor_nmos t7673(n_1591_v, n_525_v, n_696_v, n_525_port_7, n_696_port_1);
  wire [`W-1:0] temp_12479;
  spice_transistor_nmos t7678(n_2093_v, a(n_2067_v), n_804_v, temp_12479, n_804_port_1);
  spice_transistor_nmos t7687(n_575_v, n_528_v, n_696_v, n_528_port_6, n_696_port_2);
  spice_transistor_nmos t7692(n_1799_v, n_953_v, reg_pch4_v, n_953_port_3, reg_pch4_port_2);
  spice_transistor_nmos t7693(n_1800_v, reg_i4_v, n_953_v, reg_i4_port_2, n_953_port_4);
  spice_transistor_nmos t7694(n_654_v, n_949_v, reg_w4_v, n_949_port_4, reg_w4_port_2);
  spice_transistor_nmos t7695(n_657_v, reg_sph4_v, n_949_v, reg_sph4_port_2, n_949_port_5);
  spice_transistor_nmos t7696(n_658_v, n_949_v, reg_iyh4_v, n_949_port_6, reg_iyh4_port_2);
  spice_transistor_nmos t7697(n_661_v, reg_ixh4_v, n_949_v, reg_ixh4_port_2, n_949_port_7);
  spice_transistor_nmos t7698(n_662_v, n_949_v, reg_d4_v, n_949_port_8, reg_d4_port_2);
  spice_transistor_nmos t7699(n_665_v, reg_dd4_v, n_949_v, reg_dd4_port_2, n_949_port_9);
  spice_transistor_nmos t7700(n_666_v, n_949_v, reg_h4_v, n_949_port_10, reg_h4_port_2);
  spice_transistor_nmos t7701(n_669_v, reg_hh4_v, n_949_v, reg_hh4_port_2, n_949_port_11);
  spice_transistor_nmos t7702(n_670_v, n_949_v, reg_b4_v, n_949_port_12, reg_b4_port_2);
  spice_transistor_nmos t7703(n_673_v, reg_bb4_v, n_949_v, reg_bb4_port_2, n_949_port_13);
  spice_transistor_nmos t7704(n_674_v, n_949_v, reg_aa4_v, n_949_port_14, reg_aa4_port_2);
  spice_transistor_nmos t7705(n_677_v, reg_a4_v, n_949_v, reg_a4_port_2, n_949_port_15);
  wire [`W-1:0] temp_12480;
  spice_transistor_nmos t7708(n_1808_v, a(n_1813_v), n_700_v, temp_12480, n_700_port_1);
  wire [`W-1:0] temp_12481;
  spice_transistor_nmos t7709(n_1793_v, n_697_v, a(n_698_v), n_697_port_4, temp_12481);
  wire [`W-1:0] temp_12482;
  wire [`W-1:0] temp_12483;
  spice_transistor_nmos t7711(n_1811_v, a(n_699_v), a(n_683_v), temp_12482, temp_12483);
  spice_transistor_nmos t7713(n_1799_v, n_703_v, n_1814_v, n_703_port_3, n_1814_port_2);
  spice_transistor_nmos t7714(n_1800_v, n_1815_v, n_703_v, n_1815_port_2, n_703_port_4);
  spice_transistor_nmos t7715(n_654_v, n_702_v, n_1816_v, n_702_port_0, n_1816_port_2);
  spice_transistor_nmos t7716(n_657_v, n_1817_v, n_702_v, n_1817_port_2, n_702_port_1);
  spice_transistor_nmos t7717(n_658_v, n_702_v, n_1818_v, n_702_port_2, n_1818_port_2);
  spice_transistor_nmos t7718(n_661_v, n_1819_v, n_702_v, n_1819_port_2, n_702_port_3);
  spice_transistor_nmos t7719(n_662_v, n_702_v, n_1820_v, n_702_port_4, n_1820_port_2);
  spice_transistor_nmos t7720(n_665_v, n_1821_v, n_702_v, n_1821_port_2, n_702_port_5);
  spice_transistor_nmos t7722(n_666_v, n_702_v, n_1822_v, n_702_port_6, n_1822_port_2);
  spice_transistor_nmos t7723(n_669_v, n_1823_v, n_702_v, n_1823_port_2, n_702_port_7);
  spice_transistor_nmos t7724(n_670_v, n_702_v, n_1824_v, n_702_port_8, n_1824_port_2);
  spice_transistor_nmos t7725(n_673_v, n_1825_v, n_702_v, n_1825_port_2, n_702_port_9);
  spice_transistor_nmos t7726(n_674_v, n_702_v, n_1826_v, n_702_port_10, n_1826_port_2);
  spice_transistor_nmos t7727(n_677_v, n_1827_v, n_702_v, n_1827_port_2, n_702_port_11);
  spice_transistor_nmos t7731(n_1785_v, n_703_v, n_702_v, n_703_port_5, n_702_port_13);
  wire [`W-1:0] temp_12484;
  spice_transistor_nmos t7732(n_2067_v, a(n_2093_v), n_804_v, temp_12484, n_804_port_2);
  wire [`W-1:0] temp_12485;
  spice_transistor_nmos t7734(n_2085_v, n_802_v, a(n_2092_v), n_802_port_3, temp_12485);
  spice_transistor_nmos t7737(n_1785_v, n_806_v, n_807_v, n_806_port_3, n_807_port_1);
  wire [`W-1:0] temp_12486;
  spice_transistor_nmos t7742(n_1812_v, n_696_v, a(n_1574_v), n_696_port_3, temp_12486);
  wire [`W-1:0] temp_12487;
  spice_transistor_nmos t7751(n_2510_v, a(n_2503_v), n_956_v, temp_12487, n_956_port_2);
  spice_transistor_nmos t7755(n_735_v, n_796_v, n_937_v, n_796_port_6, n_937_port_8);
  spice_transistor_nmos t7762(n_1785_v, n_958_v, n_959_v, n_958_port_2, n_959_port_1);
  wire [`W-1:0] temp_12488;
  spice_transistor_nmos t7769(n_1813_v, n_700_v, a(n_1808_v), n_700_port_2, temp_12488);
  spice_transistor_nmos t7771(n_1799_v, n_958_v, reg_pch5_v, n_958_port_3, reg_pch5_port_2);
  spice_transistor_nmos t7774(n_1800_v, reg_i5_v, n_958_v, reg_i5_port_2, n_958_port_4);
  wire [`W-1:0] temp_12489;
  spice_transistor_nmos t7778(n_712_v, a(n_759_v), n_701_v, temp_12489, n_701_port_2);
  spice_transistor_nmos t7780(n_1799_v, n_806_v, n_2094_v, n_806_port_4, n_2094_port_2);
  spice_transistor_nmos t7781(n_654_v, n_959_v, reg_w5_v, n_959_port_4, reg_w5_port_2);
  spice_transistor_nmos t7782(n_1800_v, n_2095_v, n_806_v, n_2095_port_2, n_806_port_5);
  spice_transistor_nmos t7784(n_657_v, reg_sph5_v, n_959_v, reg_sph5_port_2, n_959_port_5);
  spice_transistor_nmos t7785(n_658_v, n_959_v, reg_iyh5_v, n_959_port_6, reg_iyh5_port_2);
  spice_transistor_nmos t7786(n_654_v, n_807_v, n_2096_v, n_807_port_3, n_2096_port_2);
  spice_transistor_nmos t7787(n_657_v, n_2097_v, n_807_v, n_2097_port_2, n_807_port_4);
  spice_transistor_nmos t7788(n_661_v, reg_ixh5_v, n_959_v, reg_ixh5_port_2, n_959_port_7);
  spice_transistor_nmos t7789(n_662_v, n_959_v, reg_d5_v, n_959_port_8, reg_d5_port_2);
  spice_transistor_nmos t7790(n_658_v, n_807_v, n_2098_v, n_807_port_5, n_2098_port_2);
  spice_transistor_nmos t7791(n_661_v, n_2099_v, n_807_v, n_2099_port_2, n_807_port_6);
  spice_transistor_nmos t7792(n_665_v, reg_dd5_v, n_959_v, reg_dd5_port_2, n_959_port_9);
  spice_transistor_nmos t7793(n_666_v, n_959_v, reg_h5_v, n_959_port_10, reg_h5_port_2);
  spice_transistor_nmos t7794(n_662_v, n_807_v, n_2100_v, n_807_port_7, n_2100_port_2);
  spice_transistor_nmos t7795(n_665_v, n_2101_v, n_807_v, n_2101_port_2, n_807_port_8);
  spice_transistor_nmos t7796(n_669_v, reg_hh5_v, n_959_v, reg_hh5_port_2, n_959_port_11);
  spice_transistor_nmos t7797(n_670_v, n_959_v, reg_b5_v, n_959_port_12, reg_b5_port_2);
  spice_transistor_nmos t7798(n_666_v, n_807_v, n_2102_v, n_807_port_9, n_2102_port_2);
  spice_transistor_nmos t7799(n_669_v, n_2103_v, n_807_v, n_2103_port_2, n_807_port_10);
  spice_transistor_nmos t7800(n_673_v, reg_bb5_v, n_959_v, reg_bb5_port_2, n_959_port_13);
  spice_transistor_nmos t7801(n_674_v, n_959_v, reg_aa5_v, n_959_port_14, reg_aa5_port_2);
  spice_transistor_nmos t7802(n_670_v, n_807_v, n_2104_v, n_807_port_11, n_2104_port_2);
  spice_transistor_nmos t7803(n_673_v, n_2105_v, n_807_v, n_2105_port_2, n_807_port_12);
  spice_transistor_nmos t7804(n_677_v, reg_a5_v, n_959_v, reg_a5_port_2, n_959_port_15);
  spice_transistor_nmos t7805(n_674_v, n_807_v, n_2106_v, n_807_port_13, n_2106_port_2);
  spice_transistor_nmos t7806(n_677_v, n_2107_v, n_807_v, n_2107_port_2, n_807_port_14);
  wire [`W-1:0] temp_12490;
  wire [`W-1:0] temp_12491;
  spice_transistor_nmos t7817(n_699_v, a(n_683_v), a(n_1811_v), temp_12490, temp_12491);
  spice_transistor_nmos t7822(n_575_v, n_701_v, n_716_v, n_701_port_3, n_716_port_7);
  wire [`W-1:0] temp_12492;
  spice_transistor_nmos t7823(n_1837_v, a(n_1832_v), n_707_v, temp_12492, n_707_port_0);
  wire [`W-1:0] temp_12493;
  spice_transistor_nmos t7828(n_2503_v, n_956_v, a(n_2510_v), n_956_port_3, temp_12493);
  spice_transistor_nmos t7829(n_643_v, n_937_v, n_772_v, n_937_port_9, n_772_port_7);
  wire [`W-1:0] temp_12494;
  spice_transistor_nmos t7833(n_2537_v, a(n_2529_v), n_963_v, temp_12494, n_963_port_2);
  spice_transistor_nmos t7834(n_750_v, n_790_v, n_808_v, n_790_port_5, n_808_port_6);
  wire [`W-1:0] temp_12495;
  spice_transistor_nmos t7835(n_1840_v, a(n_1835_v), n_709_v, temp_12495, n_709_port_3);
  spice_transistor_nmos t7838(n_1799_v, n_810_v, n_2119_v, n_810_port_3, n_2119_port_2);
  spice_transistor_nmos t7839(n_1800_v, n_2120_v, n_810_v, n_2120_port_2, n_810_port_4);
  spice_transistor_nmos t7840(n_654_v, n_809_v, n_2121_v, n_809_port_0, n_2121_port_2);
  spice_transistor_nmos t7841(n_657_v, n_2122_v, n_809_v, n_2122_port_2, n_809_port_1);
  spice_transistor_nmos t7842(n_658_v, n_809_v, n_2123_v, n_809_port_2, n_2123_port_2);
  spice_transistor_nmos t7843(n_661_v, n_2124_v, n_809_v, n_2124_port_2, n_809_port_3);
  spice_transistor_nmos t7844(n_662_v, n_809_v, n_2125_v, n_809_port_4, n_2125_port_2);
  spice_transistor_nmos t7845(n_665_v, n_2126_v, n_809_v, n_2126_port_2, n_809_port_5);
  spice_transistor_nmos t7846(n_666_v, n_809_v, n_2127_v, n_809_port_6, n_2127_port_2);
  spice_transistor_nmos t7847(n_669_v, n_2128_v, n_809_v, n_2128_port_2, n_809_port_7);
  spice_transistor_nmos t7848(n_670_v, n_809_v, n_2129_v, n_809_port_8, n_2129_port_2);
  spice_transistor_nmos t7849(n_673_v, n_2130_v, n_809_v, n_2130_port_2, n_809_port_9);
  spice_transistor_nmos t7850(n_674_v, n_809_v, n_2131_v, n_809_port_10, n_2131_port_2);
  spice_transistor_nmos t7851(n_677_v, n_2132_v, n_809_v, n_2132_port_2, n_809_port_11);
  wire [`W-1:0] temp_12496;
  spice_transistor_nmos t7852(n_2538_v, a(n_2512_v), n_964_v, temp_12496, n_964_port_1);
  spice_transistor_nmos t7854(n_1785_v, n_810_v, n_809_v, n_810_port_5, n_809_port_13);
  wire [`W-1:0] temp_12497;
  spice_transistor_nmos t7858(v(clk_v), n_696_v, a(n_1862_v), n_696_port_4, temp_12497);
  wire [`W-1:0] temp_12498;
  spice_transistor_nmos t7862(v(clk_v), n_701_v, a(n_737_v), n_701_port_4, temp_12498);
  wire [`W-1:0] temp_12499;
  spice_transistor_nmos t7871(n_1639_v, a(n_569_v), n_1590_v, temp_12499, n_1590_port_1);
  wire [`W-1:0] temp_12500;
  spice_transistor_nmos t7872(n_569_v, n_1590_v, a(n_1639_v), n_1590_port_2, temp_12500);
  wire [`W-1:0] temp_12501;
  spice_transistor_nmos t7885(v(clk_v), n_697_v, a(n_1858_v), n_697_port_5, temp_12501);
  wire [`W-1:0] temp_12502;
  spice_transistor_nmos t7890(n_2512_v, a(n_2538_v), n_964_v, temp_12502, n_964_port_2);
  wire [`W-1:0] temp_12503;
  spice_transistor_nmos t7892(n_2139_v, a(n_2135_v), n_833_v, temp_12503, n_833_port_0);
  wire [`W-1:0] temp_12504;
  spice_transistor_nmos t7894(n_2529_v, n_963_v, a(n_2537_v), n_963_port_3, temp_12504);
  spice_transistor_nmos t7900(n_1785_v, n_969_v, n_970_v, n_969_port_3, n_970_port_1);
  wire [`W-1:0] temp_12505;
  spice_transistor_nmos t7904(n_2141_v, a(n_2138_v), n_835_v, temp_12505, n_835_port_1);
  spice_transistor_nmos t7912(n_643_v, n_808_v, n_951_v, n_808_port_7, n_951_port_2);
  wire [`W-1:0] temp_12506;
  spice_transistor_nmos t7922(n_1835_v, a(n_1840_v), n_709_v, temp_12506, n_709_port_4);
  spice_transistor_nmos t7932(n_1785_v, n_713_v, n_708_v, n_713_port_1, n_708_port_1);
  wire [`W-1:0] temp_12507;
  spice_transistor_nmos t7937(n_680_v, a(n_1829_v), n_689_v, temp_12507, n_689_port_4);
  wire [`W-1:0] temp_12508;
  spice_transistor_nmos t7939(n_1832_v, n_707_v, a(n_1837_v), n_707_port_1, temp_12508);
  spice_transistor_nmos t7943(n_1799_v, n_969_v, n_2539_v, n_969_port_4, n_2539_port_2);
  spice_transistor_nmos t7944(n_1800_v, n_2540_v, n_969_v, n_2540_port_2, n_969_port_5);
  spice_transistor_nmos t7947(n_654_v, n_970_v, n_2541_v, n_970_port_3, n_2541_port_2);
  spice_transistor_nmos t7948(n_657_v, n_2542_v, n_970_v, n_2542_port_2, n_970_port_4);
  spice_transistor_nmos t7949(n_658_v, n_970_v, n_2543_v, n_970_port_5, n_2543_port_2);
  spice_transistor_nmos t7950(n_661_v, n_2544_v, n_970_v, n_2544_port_2, n_970_port_6);
  spice_transistor_nmos t7951(n_662_v, n_970_v, n_2545_v, n_970_port_7, n_2545_port_2);
  spice_transistor_nmos t7952(n_665_v, n_2546_v, n_970_v, n_2546_port_2, n_970_port_8);
  spice_transistor_nmos t7953(n_666_v, n_970_v, n_2547_v, n_970_port_9, n_2547_port_2);
  spice_transistor_nmos t7954(n_669_v, n_2548_v, n_970_v, n_2548_port_2, n_970_port_10);
  spice_transistor_nmos t7955(n_670_v, n_970_v, n_2549_v, n_970_port_11, n_2549_port_2);
  spice_transistor_nmos t7956(n_673_v, n_2550_v, n_970_v, n_2550_port_2, n_970_port_12);
  spice_transistor_nmos t7957(n_674_v, n_970_v, n_2551_v, n_970_port_13, n_2551_port_2);
  spice_transistor_nmos t7958(n_677_v, n_2552_v, n_970_v, n_2552_port_2, n_970_port_14);
  spice_transistor_nmos t7963(n_735_v, n_951_v, n_839_v, n_951_port_3, n_839_port_5);
  wire [`W-1:0] temp_12509;
  spice_transistor_nmos t7967(n_2138_v, a(n_2141_v), n_835_v, temp_12509, n_835_port_2);
  spice_transistor_nmos t7969(n_750_v, n_716_v, n_836_v, n_716_port_8, n_836_port_6);
  spice_transistor_nmos t7973(n_1799_v, n_713_v, reg_pcl0_v, n_713_port_3, reg_pcl0_port_2);
  spice_transistor_nmos t7974(n_1800_v, reg_r0_v, n_713_v, reg_r0_port_2, n_713_port_4);
  spice_transistor_nmos t7975(n_654_v, n_708_v, reg_z0_v, n_708_port_4, reg_z0_port_2);
  spice_transistor_nmos t7976(n_1785_v, n_841_v, n_834_v, n_841_port_1, n_834_port_1);
  wire [`W-1:0] temp_12510;
  spice_transistor_nmos t7978(n_2135_v, n_833_v, a(n_2139_v), n_833_port_1, temp_12510);
  spice_transistor_nmos t7979(n_657_v, reg_spl0_v, n_708_v, reg_spl0_port_2, n_708_port_5);
  spice_transistor_nmos t7981(n_658_v, n_708_v, reg_iyl0_v, n_708_port_6, reg_iyl0_port_2);
  spice_transistor_nmos t7982(n_661_v, reg_ixl0_v, n_708_v, reg_ixl0_port_2, n_708_port_7);
  spice_transistor_nmos t7983(n_662_v, n_708_v, reg_e0_v, n_708_port_8, reg_e0_port_2);
  spice_transistor_nmos t7985(n_665_v, reg_ee0_v, n_708_v, reg_ee0_port_2, n_708_port_9);
  spice_transistor_nmos t7986(n_666_v, n_708_v, reg_l0_v, n_708_port_10, reg_l0_port_2);
  spice_transistor_nmos t7987(n_669_v, reg_ll0_v, n_708_v, reg_ll0_port_2, n_708_port_11);
  spice_transistor_nmos t7988(n_670_v, n_708_v, reg_c0_v, n_708_port_12, reg_c0_port_2);
  spice_transistor_nmos t7989(n_673_v, reg_cc0_v, n_708_v, reg_cc0_port_2, n_708_port_13);
  spice_transistor_nmos t7991(n_674_v, n_708_v, reg_ff0_v, n_708_port_14, reg_ff0_port_2);
  spice_transistor_nmos t7992(n_734_v, n_525_v, n_837_v, n_525_port_8, n_837_port_1);
  spice_transistor_nmos t7993(n_677_v, reg_f0_v, n_708_v, reg_f0_port_2, n_708_port_15);
  spice_transistor_nmos t7997(n_1799_v, n_841_v, reg_pcl6_v, n_841_port_3, reg_pcl6_port_2);
  spice_transistor_nmos t7999(n_1799_v, n_974_v, n_2573_v, n_974_port_3, n_2573_port_2);
  spice_transistor_nmos t8000(n_1800_v, n_2574_v, n_974_v, n_2574_port_2, n_974_port_4);
  spice_transistor_nmos t8001(n_654_v, n_973_v, n_2575_v, n_973_port_0, n_2575_port_2);
  spice_transistor_nmos t8002(n_657_v, n_2576_v, n_973_v, n_2576_port_2, n_973_port_1);
  spice_transistor_nmos t8003(n_658_v, n_973_v, n_2577_v, n_973_port_2, n_2577_port_2);
  spice_transistor_nmos t8004(n_661_v, n_2578_v, n_973_v, n_2578_port_2, n_973_port_3);
  spice_transistor_nmos t8005(n_662_v, n_973_v, n_2579_v, n_973_port_4, n_2579_port_2);
  spice_transistor_nmos t8006(n_665_v, n_2580_v, n_973_v, n_2580_port_2, n_973_port_5);
  spice_transistor_nmos t8007(n_666_v, n_973_v, n_2581_v, n_973_port_6, n_2581_port_2);
  spice_transistor_nmos t8008(n_669_v, n_2582_v, n_973_v, n_2582_port_2, n_973_port_7);
  spice_transistor_nmos t8009(n_670_v, n_973_v, n_2583_v, n_973_port_8, n_2583_port_2);
  spice_transistor_nmos t8010(n_673_v, n_2584_v, n_973_v, n_2584_port_2, n_973_port_9);
  spice_transistor_nmos t8011(n_674_v, n_973_v, n_2585_v, n_973_port_10, n_2585_port_2);
  spice_transistor_nmos t8012(n_677_v, n_2586_v, n_973_v, n_2586_port_2, n_973_port_11);
  spice_transistor_nmos t8014(n_1800_v, reg_r6_v, n_841_v, reg_r6_port_2, n_841_port_4);
  spice_transistor_nmos t8015(n_654_v, n_834_v, reg_z6_v, n_834_port_4, reg_z6_port_2);
  spice_transistor_nmos t8016(n_657_v, reg_spl6_v, n_834_v, reg_spl6_port_2, n_834_port_5);
  spice_transistor_nmos t8017(n_658_v, n_834_v, reg_iyl6_v, n_834_port_6, reg_iyl6_port_2);
  spice_transistor_nmos t8018(n_1785_v, n_974_v, n_973_v, n_974_port_5, n_973_port_13);
  spice_transistor_nmos t8020(n_661_v, reg_ixl6_v, n_834_v, reg_ixl6_port_2, n_834_port_7);
  spice_transistor_nmos t8021(n_662_v, n_834_v, reg_e6_v, n_834_port_8, reg_e6_port_2);
  spice_transistor_nmos t8022(n_665_v, reg_ee6_v, n_834_v, reg_ee6_port_2, n_834_port_9);
  spice_transistor_nmos t8023(n_666_v, n_834_v, reg_l6_v, n_834_port_10, reg_l6_port_2);
  spice_transistor_nmos t8024(n_669_v, reg_ll6_v, n_834_v, reg_ll6_port_2, n_834_port_11);
  spice_transistor_nmos t8026(n_670_v, n_834_v, reg_c6_v, n_834_port_12, reg_c6_port_2);
  spice_transistor_nmos t8027(n_673_v, reg_cc6_v, n_834_v, reg_cc6_port_2, n_834_port_13);
  spice_transistor_nmos t8028(n_674_v, n_834_v, reg_ff6_v, n_834_port_14, reg_ff6_port_2);
  spice_transistor_nmos t8029(n_677_v, reg_f6_v, n_834_v, reg_f6_port_2, n_834_port_15);
  spice_transistor_nmos t8033(n_750_v, n_839_v, n_525_v, n_839_port_6, n_525_port_9);
  wire [`W-1:0] temp_12511;
  spice_transistor_nmos t8057(n_740_v, n_845_v, a(n_843_v), n_845_port_2, temp_12511);
  wire [`W-1:0] temp_12512;
  spice_transistor_nmos t8061(n_740_v, a(n_2188_v), n_850_v, temp_12512, n_850_port_2);
  spice_transistor_nmos t8064(n_820_v, n_837_v, n_845_v, n_837_port_5, n_845_port_3);
  wire [`W-1:0] temp_12513;
  spice_transistor_nmos t8067(n_2593_v, a(n_2589_v), n_979_v, temp_12513, n_979_port_0);
  spice_transistor_nmos t8068(n_604_v, n_837_v, n_850_v, n_837_port_6, n_850_port_3);
  wire [`W-1:0] temp_12514;
  spice_transistor_nmos t8077(n_2596_v, a(n_2592_v), n_981_v, temp_12514, n_981_port_1);
  spice_transistor_nmos t8079(n_1785_v, n_846_v, n_847_v, n_846_port_2, n_847_port_1);
  wire [`W-1:0] temp_12515;
  spice_transistor_nmos t8083(v(clk_v), n_845_v, a(n_2193_v), n_845_port_4, temp_12515);
  wire [`W-1:0] temp_12516;
  spice_transistor_nmos t8084(v(clk_v), n_850_v, a(n_2192_v), n_850_port_4, temp_12516);
  spice_transistor_nmos t8086(n_1799_v, n_846_v, reg_pcl7_v, n_846_port_3, reg_pcl7_port_2);
  spice_transistor_nmos t8089(n_1800_v, reg_r7_v, n_846_v, reg_r7_port_2, n_846_port_4);
  spice_transistor_nmos t8096(n_654_v, n_847_v, reg_z7_v, n_847_port_4, reg_z7_port_2);
  spice_transistor_nmos t8098(n_793_v, n_836_v, n_951_v, n_836_port_7, n_951_port_5);
  spice_transistor_nmos t8103(n_657_v, reg_spl7_v, n_847_v, reg_spl7_port_2, n_847_port_5);
  spice_transistor_nmos t8104(n_658_v, n_847_v, reg_iyl7_v, n_847_port_6, reg_iyl7_port_2);
  spice_transistor_nmos t8108(n_661_v, reg_ixl7_v, n_847_v, reg_ixl7_port_2, n_847_port_7);
  spice_transistor_nmos t8109(n_662_v, n_847_v, reg_e7_v, n_847_port_8, reg_e7_port_2);
  spice_transistor_nmos t8112(n_665_v, reg_ee7_v, n_847_v, reg_ee7_port_2, n_847_port_9);
  spice_transistor_nmos t8113(n_666_v, n_847_v, reg_l7_v, n_847_port_10, reg_l7_port_2);
  spice_transistor_nmos t8114(n_1785_v, n_714_v, n_715_v, n_714_port_2, n_715_port_1);
  spice_transistor_nmos t8116(n_669_v, reg_ll7_v, n_847_v, reg_ll7_port_2, n_847_port_11);
  spice_transistor_nmos t8117(n_670_v, n_847_v, reg_c7_v, n_847_port_12, reg_c7_port_2);
  spice_transistor_nmos t8120(n_673_v, reg_cc7_v, n_847_v, reg_cc7_port_2, n_847_port_13);
  wire [`W-1:0] temp_12517;
  spice_transistor_nmos t8121(v(clk_v), a(n_2567_v), n_966_v, temp_12517, n_966_port_2);
  spice_transistor_nmos t8122(n_674_v, n_847_v, reg_ff7_v, n_847_port_14, reg_ff7_port_2);
  spice_transistor_nmos t8125(n_677_v, reg_f7_v, n_847_v, reg_f7_port_2, n_847_port_15);
  spice_transistor_nmos t8127(n_1799_v, n_714_v, reg_pcl1_v, n_714_port_3, reg_pcl1_port_2);
  spice_transistor_nmos t8133(n_1800_v, reg_r1_v, n_714_v, reg_r1_port_2, n_714_port_4);
  wire [`W-1:0] temp_12518;
  spice_transistor_nmos t8135(n_740_v, a(n_2570_v), n_966_v, temp_12518, n_966_port_3);
  spice_transistor_nmos t8136(n_793_v, n_837_v, n_755_v, n_837_port_8, n_755_port_6);
  spice_transistor_nmos t8137(n_820_v, n_966_v, n_951_v, n_966_port_4, n_951_port_8);
  wire [`W-1:0] temp_12519;
  spice_transistor_nmos t8139(n_2592_v, a(n_2596_v), n_981_v, temp_12519, n_981_port_2);
  spice_transistor_nmos t8140(n_646_v, n_2504_v, n_951_v, n_2504_port_5, n_951_port_10);
  spice_transistor_nmos t8146(n_654_v, n_715_v, reg_z1_v, n_715_port_4, reg_z1_port_2);
  spice_transistor_nmos t8147(n_1785_v, n_982_v, n_980_v, n_982_port_1, n_980_port_1);
  wire [`W-1:0] temp_12520;
  spice_transistor_nmos t8149(n_2589_v, n_979_v, a(n_2593_v), n_979_port_1, temp_12520);
  spice_transistor_nmos t8152(n_657_v, reg_spl1_v, n_715_v, reg_spl1_port_2, n_715_port_5);
  spice_transistor_nmos t8156(n_658_v, n_715_v, reg_iyl1_v, n_715_port_6, reg_iyl1_port_2);
  wire [`W-1:0] temp_12521;
  spice_transistor_nmos t8159(n_2194_v, a(n_2180_v), n_856_v, temp_12521, n_856_port_3);
  spice_transistor_nmos t8160(n_661_v, reg_ixl1_v, n_715_v, reg_ixl1_port_2, n_715_port_7);
  spice_transistor_nmos t8162(n_662_v, n_715_v, reg_e1_v, n_715_port_8, reg_e1_port_2);
  spice_transistor_nmos t8166(n_1799_v, n_982_v, reg_pch6_v, n_982_port_3, reg_pch6_port_2);
  spice_transistor_nmos t8167(n_1800_v, reg_i6_v, n_982_v, reg_i6_port_2, n_982_port_4);
  spice_transistor_nmos t8168(n_654_v, n_980_v, reg_w6_v, n_980_port_4, reg_w6_port_2);
  spice_transistor_nmos t8169(n_657_v, reg_sph6_v, n_980_v, reg_sph6_port_2, n_980_port_5);
  spice_transistor_nmos t8170(n_658_v, n_980_v, reg_iyh6_v, n_980_port_6, reg_iyh6_port_2);
  spice_transistor_nmos t8171(n_661_v, reg_ixh6_v, n_980_v, reg_ixh6_port_2, n_980_port_7);
  spice_transistor_nmos t8172(n_662_v, n_980_v, reg_d6_v, n_980_port_8, reg_d6_port_2);
  spice_transistor_nmos t8173(n_665_v, reg_dd6_v, n_980_v, reg_dd6_port_2, n_980_port_9);
  spice_transistor_nmos t8174(n_666_v, n_980_v, reg_h6_v, n_980_port_10, reg_h6_port_2);
  spice_transistor_nmos t8175(n_669_v, reg_hh6_v, n_980_v, reg_hh6_port_2, n_980_port_11);
  spice_transistor_nmos t8176(n_670_v, n_980_v, reg_b6_v, n_980_port_12, reg_b6_port_2);
  spice_transistor_nmos t8177(n_673_v, reg_bb6_v, n_980_v, reg_bb6_port_2, n_980_port_13);
  spice_transistor_nmos t8178(n_674_v, n_980_v, reg_aa6_v, n_980_port_14, reg_aa6_port_2);
  spice_transistor_nmos t8179(n_677_v, reg_a6_v, n_980_v, reg_a6_port_2, n_980_port_15);
  spice_transistor_nmos t8181(n_665_v, reg_ee1_v, n_715_v, reg_ee1_port_2, n_715_port_9);
  spice_transistor_nmos t8182(n_666_v, n_715_v, reg_l1_v, n_715_port_10, reg_l1_port_2);
  spice_transistor_nmos t8185(n_669_v, reg_ll1_v, n_715_v, reg_ll1_port_2, n_715_port_11);
  spice_transistor_nmos t8186(n_670_v, n_715_v, reg_c1_v, n_715_port_12, reg_c1_port_2);
  spice_transistor_nmos t8189(n_673_v, reg_cc1_v, n_715_v, reg_cc1_port_2, n_715_port_13);
  spice_transistor_nmos t8190(n_674_v, n_715_v, reg_ff1_v, n_715_port_14, reg_ff1_port_2);
  spice_transistor_nmos t8193(n_677_v, reg_f1_v, n_715_v, reg_f1_port_2, n_715_port_15);
  wire [`W-1:0] temp_12522;
  spice_transistor_nmos t8201(n_2195_v, a(n_2164_v), n_857_v, temp_12522, n_857_port_1);
  spice_transistor_nmos t8212(n_1785_v, n_984_v, n_985_v, n_984_port_2, n_985_port_1);
  spice_transistor_nmos t8218(n_1799_v, n_984_v, reg_pch7_v, n_984_port_3, reg_pch7_port_2);
  wire [`W-1:0] temp_12523;
  spice_transistor_nmos t8220(n_1888_v, a(n_1865_v), n_721_v, temp_12523, n_721_port_2);
  spice_transistor_nmos t8221(n_1800_v, reg_i7_v, n_984_v, reg_i7_port_2, n_984_port_4);
  spice_transistor_nmos t8225(n_654_v, n_985_v, reg_w7_v, n_985_port_4, reg_w7_port_2);
  spice_transistor_nmos t8228(n_657_v, reg_sph7_v, n_985_v, reg_sph7_port_2, n_985_port_5);
  spice_transistor_nmos t8229(n_658_v, n_985_v, reg_iyh7_v, n_985_port_6, reg_iyh7_port_2);
  spice_transistor_nmos t8232(n_661_v, reg_ixh7_v, n_985_v, reg_ixh7_port_2, n_985_port_7);
  spice_transistor_nmos t8233(n_662_v, n_985_v, reg_d7_v, n_985_port_8, reg_d7_port_2);
  spice_transistor_nmos t8236(n_665_v, reg_dd7_v, n_985_v, reg_dd7_port_2, n_985_port_9);
  spice_transistor_nmos t8237(n_666_v, n_985_v, reg_h7_v, n_985_port_10, reg_h7_port_2);
  spice_transistor_nmos t8240(n_669_v, reg_hh7_v, n_985_v, reg_hh7_port_2, n_985_port_11);
  spice_transistor_nmos t8241(n_670_v, n_985_v, reg_b7_v, n_985_port_12, reg_b7_port_2);
  spice_transistor_nmos t8244(n_673_v, reg_bb7_v, n_985_v, reg_bb7_port_2, n_985_port_13);
  spice_transistor_nmos t8245(n_674_v, n_985_v, reg_aa7_v, n_985_port_14, reg_aa7_port_2);
  spice_transistor_nmos t8248(n_677_v, reg_a7_v, n_985_v, reg_a7_port_2, n_985_port_15);
  wire [`W-1:0] temp_12524;
  spice_transistor_nmos t8255(n_1889_v, a(n_1866_v), n_722_v, temp_12524, n_722_port_1);
  wire [`W-1:0] temp_12525;
  spice_transistor_nmos t8256(n_740_v, n_988_v, a(n_986_v), n_988_port_1, temp_12525);
  wire [`W-1:0] temp_12526;
  spice_transistor_nmos t8261(n_740_v, a(n_2661_v), n_993_v, temp_12526, n_993_port_2);
  spice_transistor_nmos t8265(n_820_v, n_983_v, n_988_v, n_983_port_4, n_988_port_2);
  spice_transistor_nmos t8268(n_604_v, n_983_v, n_993_v, n_983_port_5, n_993_port_3);
  wire [`W-1:0] temp_12527;
  spice_transistor_nmos t8270(n_1763_v, n_726_v, a(n_727_v), n_726_port_2, temp_12527);
  wire [`W-1:0] temp_12528;
  spice_transistor_nmos t8275(v(clk_v), n_988_v, a(n_2666_v), n_988_port_4, temp_12528);
  wire [`W-1:0] temp_12529;
  spice_transistor_nmos t8279(v(clk_v), n_993_v, a(n_2667_v), n_993_port_4, temp_12529);
  wire [`W-1:0] temp_12530;
  spice_transistor_nmos t8283(n_2164_v, a(n_2195_v), n_857_v, temp_12530, n_857_port_2);
  wire [`W-1:0] temp_12531;
  spice_transistor_nmos t8285(n_680_v, a(n_2220_v), n_2116_v, temp_12531, n_2116_port_3);
  wire [`W-1:0] temp_12532;
  spice_transistor_nmos t8286(n_2180_v, n_856_v, a(n_2194_v), n_856_port_4, temp_12532);
  wire [`W-1:0] temp_12533;
  spice_transistor_nmos t8288(n_2218_v, a(n_2213_v), n_861_v, temp_12533, n_861_port_1);
  spice_transistor_nmos t8291(n_735_v, n_772_v, n_837_v, n_772_port_8, n_837_port_9);
  spice_transistor_nmos t8293(n_1785_v, n_863_v, n_864_v, n_863_port_3, n_864_port_1);
  wire [`W-1:0] temp_12534;
  spice_transistor_nmos t8297(n_2642_v, a(n_2618_v), n_994_v, temp_12534, n_994_port_1);
  spice_transistor_nmos t8304(n_793_v, n_983_v, n_796_v, n_983_port_7, n_796_port_7);
  spice_transistor_nmos t8310(n_575_v, n_545_v, n_726_v, n_545_port_8, n_726_port_3);
  wire [`W-1:0] temp_12535;
  spice_transistor_nmos t8317(n_1794_v, a(n_765_v), n_726_v, temp_12535, n_726_port_4);
  wire [`W-1:0] temp_12536;
  spice_transistor_nmos t8319(n_680_v, n_723_v, a(n_1907_v), n_723_port_4, temp_12536);
  wire [`W-1:0] temp_12537;
  spice_transistor_nmos t8326(n_1866_v, a(n_1889_v), n_722_v, temp_12537, n_722_port_2);
  wire [`W-1:0] temp_12538;
  spice_transistor_nmos t8332(n_1904_v, a(n_1908_v), n_728_v, temp_12538, n_728_port_2);
  wire [`W-1:0] temp_12539;
  spice_transistor_nmos t8333(n_1865_v, n_721_v, a(n_1888_v), n_721_port_3, temp_12539);
  spice_transistor_nmos t8340(n_1799_v, n_863_v, n_2196_v, n_863_port_4, n_2196_port_2);
  spice_transistor_nmos t8341(n_1800_v, n_2197_v, n_863_v, n_2197_port_2, n_863_port_5);
  wire [`W-1:0] temp_12540;
  spice_transistor_nmos t8346(n_2618_v, a(n_2642_v), n_994_v, temp_12540, n_994_port_2);
  spice_transistor_nmos t8349(n_1785_v, n_731_v, n_732_v, n_731_port_3, n_732_port_1);
  spice_transistor_nmos t8350(n_654_v, n_864_v, n_2198_v, n_864_port_3, n_2198_port_2);
  spice_transistor_nmos t8352(n_657_v, n_2199_v, n_864_v, n_2199_port_2, n_864_port_4);
  spice_transistor_nmos t8353(n_658_v, n_864_v, n_2200_v, n_864_port_5, n_2200_port_2);
  spice_transistor_nmos t8354(n_1785_v, n_998_v, n_999_v, n_998_port_3, n_999_port_1);
  spice_transistor_nmos t8355(n_661_v, n_2201_v, n_864_v, n_2201_port_2, n_864_port_6);
  spice_transistor_nmos t8356(n_662_v, n_864_v, n_2202_v, n_864_port_7, n_2202_port_2);
  spice_transistor_nmos t8357(n_665_v, n_2203_v, n_864_v, n_2203_port_2, n_864_port_8);
  spice_transistor_nmos t8358(n_666_v, n_864_v, n_2204_v, n_864_port_9, n_2204_port_2);
  spice_transistor_nmos t8359(n_669_v, n_2205_v, n_864_v, n_2205_port_2, n_864_port_10);
  spice_transistor_nmos t8360(n_670_v, n_864_v, n_2206_v, n_864_port_11, n_2206_port_2);
  spice_transistor_nmos t8361(n_673_v, n_2207_v, n_864_v, n_2207_port_2, n_864_port_12);
  spice_transistor_nmos t8362(n_674_v, n_864_v, n_2208_v, n_864_port_13, n_2208_port_2);
  spice_transistor_nmos t8363(n_677_v, n_2209_v, n_864_v, n_2209_port_2, n_864_port_14);
  wire [`W-1:0] temp_12541;
  spice_transistor_nmos t8371(n_2213_v, n_861_v, a(n_2218_v), n_861_port_2, temp_12541);
  wire [`W-1:0] temp_12542;
  spice_transistor_nmos t8386(n_2675_v, a(n_2670_v), n_1001_v, temp_12542, n_1001_port_2);
  spice_transistor_nmos t8390(n_735_v, n_803_v, n_983_v, n_803_port_7, n_983_port_8);
  wire [`W-1:0] temp_12543;
  spice_transistor_nmos t8395(n_1908_v, n_728_v, a(n_1904_v), n_728_port_3, temp_12543);
  spice_transistor_nmos t8398(n_1799_v, n_998_v, n_2643_v, n_998_port_4, n_2643_port_2);
  spice_transistor_nmos t8399(n_1800_v, n_2644_v, n_998_v, n_2644_port_2, n_998_port_5);
  spice_transistor_nmos t8401(n_654_v, n_999_v, n_2645_v, n_999_port_3, n_2645_port_2);
  spice_transistor_nmos t8402(n_657_v, n_2646_v, n_999_v, n_2646_port_2, n_999_port_4);
  spice_transistor_nmos t8403(n_658_v, n_999_v, n_2647_v, n_999_port_5, n_2647_port_2);
  spice_transistor_nmos t8404(n_661_v, n_2648_v, n_999_v, n_2648_port_2, n_999_port_6);
  spice_transistor_nmos t8405(n_662_v, n_999_v, n_2649_v, n_999_port_7, n_2649_port_2);
  spice_transistor_nmos t8406(n_665_v, n_2650_v, n_999_v, n_2650_port_2, n_999_port_8);
  spice_transistor_nmos t8407(n_666_v, n_999_v, n_2651_v, n_999_port_9, n_2651_port_2);
  spice_transistor_nmos t8408(n_669_v, n_2652_v, n_999_v, n_2652_port_2, n_999_port_10);
  spice_transistor_nmos t8409(n_670_v, n_999_v, n_2653_v, n_999_port_11, n_2653_port_2);
  spice_transistor_nmos t8410(n_673_v, n_2654_v, n_999_v, n_2654_port_2, n_999_port_12);
  spice_transistor_nmos t8411(n_674_v, n_999_v, n_2655_v, n_999_port_13, n_2655_port_2);
  spice_transistor_nmos t8412(n_677_v, n_2656_v, n_999_v, n_2656_port_2, n_999_port_14);
  spice_transistor_nmos t8422(n_1799_v, n_731_v, n_1890_v, n_731_port_4, n_1890_port_2);
  spice_transistor_nmos t8423(n_1800_v, n_1891_v, n_731_v, n_1891_port_2, n_731_port_5);
  spice_transistor_nmos t8425(n_643_v, n_796_v, n_852_v, n_796_port_8, n_852_port_2);
  spice_transistor_nmos t8428(n_654_v, n_732_v, n_1892_v, n_732_port_3, n_1892_port_2);
  spice_transistor_nmos t8432(n_657_v, n_1893_v, n_732_v, n_1893_port_2, n_732_port_4);
  spice_transistor_nmos t8434(n_658_v, n_732_v, n_1894_v, n_732_port_5, n_1894_port_2);
  spice_transistor_nmos t8435(n_661_v, n_1895_v, n_732_v, n_1895_port_2, n_732_port_6);
  spice_transistor_nmos t8436(n_662_v, n_732_v, n_1896_v, n_732_port_7, n_1896_port_2);
  spice_transistor_nmos t8437(n_643_v, n_983_v, n_783_v, n_983_port_9, n_783_port_8);
  spice_transistor_nmos t8438(n_665_v, n_1897_v, n_732_v, n_1897_port_2, n_732_port_8);
  spice_transistor_nmos t8439(n_666_v, n_732_v, n_1898_v, n_732_port_9, n_1898_port_2);
  spice_transistor_nmos t8441(n_669_v, n_1899_v, n_732_v, n_1899_port_2, n_732_port_10);
  spice_transistor_nmos t8442(n_670_v, n_732_v, n_1900_v, n_732_port_11, n_1900_port_2);
  spice_transistor_nmos t8444(n_673_v, n_1901_v, n_732_v, n_1901_port_2, n_732_port_12);
  spice_transistor_nmos t8445(n_674_v, n_732_v, n_1902_v, n_732_port_13, n_1902_port_2);
  spice_transistor_nmos t8449(n_677_v, n_1903_v, n_732_v, n_1903_port_2, n_732_port_14);
  wire [`W-1:0] temp_12544;
  spice_transistor_nmos t8451(n_2670_v, n_1001_v, a(n_2675_v), n_1001_port_3, temp_12544);
  spice_transistor_nmos t8454(n_1799_v, n_871_v, n_2232_v, n_871_port_3, n_2232_port_2);
  spice_transistor_nmos t8455(n_1800_v, n_2233_v, n_871_v, n_2233_port_2, n_871_port_4);
  spice_transistor_nmos t8456(n_654_v, n_870_v, n_2234_v, n_870_port_0, n_2234_port_2);
  spice_transistor_nmos t8457(n_657_v, n_2235_v, n_870_v, n_2235_port_2, n_870_port_1);
  spice_transistor_nmos t8458(n_658_v, n_870_v, n_2236_v, n_870_port_2, n_2236_port_2);
  spice_transistor_nmos t8460(n_661_v, n_2237_v, n_870_v, n_2237_port_2, n_870_port_3);
  spice_transistor_nmos t8461(n_662_v, n_870_v, n_2238_v, n_870_port_4, n_2238_port_2);
  spice_transistor_nmos t8462(n_665_v, n_2239_v, n_870_v, n_2239_port_2, n_870_port_5);
  spice_transistor_nmos t8463(n_666_v, n_870_v, n_2240_v, n_870_port_6, n_2240_port_2);
  spice_transistor_nmos t8464(n_669_v, n_2241_v, n_870_v, n_2241_port_2, n_870_port_7);
  spice_transistor_nmos t8465(n_643_v, n_995_v, n_836_v, n_995_port_2, n_836_port_8);
  spice_transistor_nmos t8466(n_670_v, n_870_v, n_2242_v, n_870_port_8, n_2242_port_2);
  spice_transistor_nmos t8467(n_673_v, n_2243_v, n_870_v, n_2243_port_2, n_870_port_9);
  spice_transistor_nmos t8468(n_674_v, n_870_v, n_2244_v, n_870_port_10, n_2244_port_2);
  spice_transistor_nmos t8469(n_677_v, n_2245_v, n_870_v, n_2245_port_2, n_870_port_11);
  spice_transistor_nmos t8470(n_793_v, n_995_v, n_839_v, n_995_port_3, n_839_port_7);
  spice_transistor_nmos t8476(n_1785_v, n_871_v, n_870_v, n_871_port_5, n_870_port_13);
  wire [`W-1:0] temp_12545;
  spice_transistor_nmos t8499(v(clk_v), n_726_v, a(n_1943_v), n_726_port_5, temp_12545);
  spice_transistor_nmos t8503(n_735_v, n_852_v, n_808_v, n_852_port_3, n_808_port_8);
  wire [`W-1:0] temp_12546;
  spice_transistor_nmos t8508(n_680_v, a(n_2689_v), n_2617_v, temp_12546, n_2617_port_4);
  spice_transistor_nmos t8518(n_1799_v, n_739_v, n_1915_v, n_739_port_3, n_1915_port_2);
  spice_transistor_nmos t8519(n_1800_v, n_1916_v, n_739_v, n_1916_port_2, n_739_port_4);
  spice_transistor_nmos t8520(n_654_v, n_738_v, n_1917_v, n_738_port_0, n_1917_port_2);
  spice_transistor_nmos t8521(n_657_v, n_1918_v, n_738_v, n_1918_port_2, n_738_port_1);
  spice_transistor_nmos t8522(n_658_v, n_738_v, n_1919_v, n_738_port_2, n_1919_port_2);
  spice_transistor_nmos t8523(n_661_v, n_1920_v, n_738_v, n_1920_port_2, n_738_port_3);
  spice_transistor_nmos t8524(n_662_v, n_738_v, n_1921_v, n_738_port_4, n_1921_port_2);
  spice_transistor_nmos t8525(n_665_v, n_1922_v, n_738_v, n_1922_port_2, n_738_port_5);
  wire [`W-1:0] temp_12547;
  spice_transistor_nmos t8527(n_2253_v, a(n_2249_v), n_879_v, temp_12547, n_879_port_0);
  spice_transistor_nmos t8528(n_666_v, n_738_v, n_1923_v, n_738_port_6, n_1923_port_2);
  spice_transistor_nmos t8529(n_669_v, n_1924_v, n_738_v, n_1924_port_2, n_738_port_7);
  spice_transistor_nmos t8530(n_670_v, n_738_v, n_1925_v, n_738_port_8, n_1925_port_2);
  spice_transistor_nmos t8531(n_673_v, n_1926_v, n_738_v, n_1926_port_2, n_738_port_9);
  spice_transistor_nmos t8532(n_735_v, n_681_v, n_995_v, n_681_port_5, n_995_port_4);
  spice_transistor_nmos t8533(n_674_v, n_738_v, n_1927_v, n_738_port_10, n_1927_port_2);
  spice_transistor_nmos t8534(n_677_v, n_1928_v, n_738_v, n_1928_port_2, n_738_port_11);
  wire [`W-1:0] temp_12548;
  spice_transistor_nmos t8537(n_2257_v, a(n_2252_v), n_881_v, temp_12548, n_881_port_2);
  spice_transistor_nmos t8543(n_1785_v, n_739_v, n_738_v, n_739_port_5, n_738_port_13);
  wire [`W-1:0] temp_12549;
  spice_transistor_nmos t8544(n_680_v, n_1009_v, a(n_2698_v), n_1009_port_4, temp_12549);
  wire [`W-1:0] temp_12550;
  spice_transistor_nmos t8545(v(clk_v), a(n_2690_v), n_1005_v, temp_12550, n_1005_port_3);
  spice_transistor_nmos t8554(n_820_v, n_1005_v, n_995_v, n_1005_port_4, n_995_port_8);
  wire [`W-1:0] temp_12551;
  spice_transistor_nmos t8555(n_740_v, a(n_2692_v), n_1005_v, temp_12551, n_1005_port_5);
  spice_transistor_nmos t8558(n_646_v, n_816_v, n_995_v, n_816_port_6, n_995_port_10);
  wire [`W-1:0] temp_12552;
  spice_transistor_nmos t8614(n_1939_v, a(n_1934_v), n_744_v, temp_12552, n_744_port_0);
  wire [`W-1:0] temp_12553;
  spice_transistor_nmos t8621(n_1941_v, a(n_1937_v), n_746_v, temp_12553, n_746_port_3);
  wire [`W-1:0] temp_12554;
  spice_transistor_nmos t8630(n_2252_v, a(n_2257_v), n_881_v, temp_12554, n_881_port_3);
  wire [`W-1:0] temp_12555;
  spice_transistor_nmos t8638(n_680_v, n_2700_v, a(n_2715_v), n_2700_port_4, temp_12555);
  spice_transistor_nmos t8641(n_1785_v, n_884_v, n_880_v, n_884_port_1, n_880_port_1);
  wire [`W-1:0] temp_12556;
  spice_transistor_nmos t8648(n_2249_v, n_879_v, a(n_2253_v), n_879_port_1, temp_12556);
  spice_transistor_nmos t8651(n_793_v, n_803_v, n_852_v, n_803_port_8, n_852_port_5);
  wire [`W-1:0] temp_12557;
  spice_transistor_nmos t8659(n_680_v, n_2701_v, a(n_2720_v), n_2701_port_4, temp_12557);
  wire [`W-1:0] temp_12558;
  spice_transistor_nmos t8660(n_680_v, n_2702_v, a(n_2721_v), n_2702_port_4, temp_12558);
  wire [`W-1:0] temp_12559;
  spice_transistor_nmos t8661(n_680_v, n_2703_v, a(n_2722_v), n_2703_port_4, temp_12559);
  wire [`W-1:0] temp_12560;
  spice_transistor_nmos t8662(n_680_v, n_2704_v, a(n_2723_v), n_2704_port_4, temp_12560);
  wire [`W-1:0] temp_12561;
  spice_transistor_nmos t8663(n_680_v, n_2705_v, a(n_2724_v), n_2705_port_4, temp_12561);
  wire [`W-1:0] temp_12562;
  spice_transistor_nmos t8664(v(clk_v), a(n_1210_v), n_181_v, temp_12562, n_181_port_6);
  spice_transistor_nmos t8672(n_1799_v, n_884_v, reg_pch0_v, n_884_port_3, reg_pch0_port_2);
  spice_transistor_nmos t8673(n_1800_v, reg_i0_v, n_884_v, reg_i0_port_2, n_884_port_4);
  spice_transistor_nmos t8674(n_654_v, n_880_v, reg_w0_v, n_880_port_4, reg_w0_port_2);
  spice_transistor_nmos t8675(n_657_v, reg_sph0_v, n_880_v, reg_sph0_port_2, n_880_port_5);
  spice_transistor_nmos t8676(n_658_v, n_880_v, reg_iyh0_v, n_880_port_6, reg_iyh0_port_2);
  spice_transistor_nmos t8677(n_661_v, reg_ixh0_v, n_880_v, reg_ixh0_port_2, n_880_port_7);
  spice_transistor_nmos t8678(n_662_v, n_880_v, reg_d0_v, n_880_port_8, reg_d0_port_2);
  spice_transistor_nmos t8679(n_665_v, reg_dd0_v, n_880_v, reg_dd0_port_2, n_880_port_9);
  spice_transistor_nmos t8680(n_666_v, n_880_v, reg_h0_v, n_880_port_10, reg_h0_port_2);
  spice_transistor_nmos t8681(n_669_v, reg_hh0_v, n_880_v, reg_hh0_port_2, n_880_port_11);
  spice_transistor_nmos t8682(n_670_v, n_880_v, reg_b0_v, n_880_port_12, reg_b0_port_2);
  spice_transistor_nmos t8683(n_673_v, reg_bb0_v, n_880_v, reg_bb0_port_2, n_880_port_13);
  spice_transistor_nmos t8684(n_674_v, n_880_v, reg_aa0_v, n_880_port_14, reg_aa0_port_2);
  spice_transistor_nmos t8685(n_677_v, reg_a0_v, n_880_v, reg_a0_port_2, n_880_port_15);
  wire [`W-1:0] temp_12563;
  spice_transistor_nmos t8691(v(clk_v), a(n_2255_v), n_867_v, temp_12563, n_867_port_1);
  wire [`W-1:0] temp_12564;
  spice_transistor_nmos t8703(n_740_v, a(n_2272_v), n_867_v, temp_12564, n_867_port_3);
  wire [`W-1:0] temp_12565;
  spice_transistor_nmos t8706(n_680_v, n_1020_v, a(n_2737_v), n_1020_port_4, temp_12565);
  wire [`W-1:0] temp_12566;
  spice_transistor_nmos t8707(n_680_v, n_1014_v, a(n_2738_v), n_1014_port_4, temp_12566);
  wire [`W-1:0] temp_12567;
  spice_transistor_nmos t8708(n_680_v, n_1017_v, a(n_2739_v), n_1017_port_4, temp_12567);
  wire [`W-1:0] temp_12568;
  spice_transistor_nmos t8709(n_680_v, n_1018_v, a(n_2740_v), n_1018_port_4, temp_12568);
  spice_transistor_nmos t8713(n_546_v, n_138_v, n_545_v, n_138_port_3, n_545_port_10);
  spice_transistor_nmos t8714(n_546_v, n_196_v, n_528_v, n_196_port_4, n_528_port_7);
  spice_transistor_nmos t8715(n_546_v, n_412_v, n_526_v, n_412_port_4, n_526_port_8);
  wire [`W-1:0] temp_12569;
  spice_transistor_nmos t8716(n_1937_v, a(n_1941_v), n_746_v, temp_12569, n_746_port_4);
  spice_transistor_nmos t8717(n_546_v, n_370_v, n_525_v, n_370_port_4, n_525_port_11);
  spice_transistor_nmos t8724(n_820_v, n_867_v, n_852_v, n_867_port_4, n_852_port_8);
  spice_transistor_nmos t8727(n_646_v, n_2211_v, n_852_v, n_2211_port_5, n_852_port_10);
  spice_transistor_nmos t8731(n_1785_v, n_749_v, n_745_v, n_749_port_1, n_745_port_1);
  spice_transistor_nmos t8732(n_1785_v, n_885_v, n_886_v, n_885_port_2, n_886_port_1);
  spice_transistor_nmos t8738(n_1799_v, n_885_v, reg_pch1_v, n_885_port_3, reg_pch1_port_2);
  spice_transistor_nmos t8741(n_1800_v, reg_i1_v, n_885_v, reg_i1_port_2, n_885_port_4);
  wire [`W-1:0] temp_12570;
  spice_transistor_nmos t8742(n_1934_v, n_744_v, a(n_1939_v), n_744_port_1, temp_12570);
  spice_transistor_nmos t8746(n_654_v, n_886_v, reg_w1_v, n_886_port_4, reg_w1_port_2);
  spice_transistor_nmos t8749(n_657_v, reg_sph1_v, n_886_v, reg_sph1_port_2, n_886_port_5);
  spice_transistor_nmos t8750(n_658_v, n_886_v, reg_iyh1_v, n_886_port_6, reg_iyh1_port_2);
  spice_transistor_nmos t8753(n_661_v, reg_ixh1_v, n_886_v, reg_ixh1_port_2, n_886_port_7);
  spice_transistor_nmos t8754(n_662_v, n_886_v, reg_d1_v, n_886_port_8, reg_d1_port_2);
  spice_transistor_nmos t8757(n_665_v, reg_dd1_v, n_886_v, reg_dd1_port_2, n_886_port_9);
  spice_transistor_nmos t8758(n_666_v, n_886_v, reg_h1_v, n_886_port_10, reg_h1_port_2);
  spice_transistor_nmos t8761(n_669_v, reg_hh1_v, n_886_v, reg_hh1_port_2, n_886_port_11);
  spice_transistor_nmos t8762(n_670_v, n_886_v, reg_b1_v, n_886_port_12, reg_b1_port_2);
  spice_transistor_nmos t8765(n_673_v, reg_bb1_v, n_886_v, reg_bb1_port_2, n_886_port_13);
  spice_transistor_nmos t8766(n_674_v, n_886_v, reg_aa1_v, n_886_port_14, reg_aa1_port_2);
  spice_transistor_nmos t8769(n_677_v, reg_a1_v, n_886_v, reg_a1_port_2, n_886_port_15);
  spice_transistor_nmos t8780(n_1799_v, n_749_v, reg_pcl2_v, n_749_port_3, reg_pcl2_port_2);
  spice_transistor_nmos t8781(n_1800_v, reg_r2_v, n_749_v, reg_r2_port_2, n_749_port_4);
  spice_transistor_nmos t8782(n_654_v, n_745_v, reg_z2_v, n_745_port_4, reg_z2_port_2);
  spice_transistor_nmos t8783(n_657_v, reg_spl2_v, n_745_v, reg_spl2_port_2, n_745_port_5);
  wire [`W-1:0] temp_12571;
  spice_transistor_nmos t8785(n_2304_v, a(n_2298_v), n_892_v, temp_12571, n_892_port_3);
  spice_transistor_nmos t8786(n_658_v, n_745_v, reg_iyl2_v, n_745_port_6, reg_iyl2_port_2);
  spice_transistor_nmos t8787(n_661_v, reg_ixl2_v, n_745_v, reg_ixl2_port_2, n_745_port_7);
  spice_transistor_nmos t8788(n_662_v, n_745_v, reg_e2_v, n_745_port_8, reg_e2_port_2);
  spice_transistor_nmos t8789(n_665_v, reg_ee2_v, n_745_v, reg_ee2_port_2, n_745_port_9);
  spice_transistor_nmos t8790(n_666_v, n_745_v, reg_l2_v, n_745_port_10, reg_l2_port_2);
  spice_transistor_nmos t8791(n_669_v, reg_ll2_v, n_745_v, reg_ll2_port_2, n_745_port_11);
  spice_transistor_nmos t8792(n_670_v, n_745_v, reg_c2_v, n_745_port_12, reg_c2_port_2);
  spice_transistor_nmos t8793(n_673_v, reg_cc2_v, n_745_v, reg_cc2_port_2, n_745_port_13);
  spice_transistor_nmos t8794(n_674_v, n_745_v, reg_ff2_v, n_745_port_14, reg_ff2_port_2);
  spice_transistor_nmos t8795(n_677_v, reg_f2_v, n_745_v, reg_f2_port_2, n_745_port_15);
  wire [`W-1:0] temp_12572;
  spice_transistor_nmos t8804(n_2305_v, a(n_2281_v), n_893_v, temp_12572, n_893_port_1);
  wire [`W-1:0] temp_12573;
  spice_transistor_nmos t8810(n_680_v, a(n_2302_v), n_2320_v, temp_12573, n_2320_port_4);
  spice_transistor_nmos t8835(n_750_v, n_545_v, n_755_v, n_545_port_11, n_755_port_7);
  wire [`W-1:0] temp_12574;
  spice_transistor_nmos t8838(n_740_v, n_897_v, a(n_894_v), n_897_port_2, temp_12574);
  wire [`W-1:0] temp_12575;
  spice_transistor_nmos t8840(n_2281_v, a(n_2305_v), n_893_v, temp_12575, n_893_port_2);
  wire [`W-1:0] temp_12576;
  spice_transistor_nmos t8842(n_740_v, a(n_2331_v), n_899_v, temp_12576, n_899_port_2);
  wire [`W-1:0] temp_12577;
  spice_transistor_nmos t8844(n_2298_v, n_892_v, a(n_2304_v), n_892_port_4, temp_12577);
  spice_transistor_nmos t8845(n_820_v, n_889_v, n_897_v, n_889_port_8, n_897_port_3);
  spice_transistor_nmos t8846(n_604_v, n_889_v, n_899_v, n_889_port_9, n_899_port_3);
  spice_transistor_nmos t8852(n_1785_v, n_901_v, n_902_v, n_901_port_5, n_902_port_13);
  spice_transistor_nmos t8855(n_1785_v, n_752_v, n_753_v, n_752_port_2, n_753_port_9);
  wire [`W-1:0] temp_12578;
  spice_transistor_nmos t8861(v(clk_v), n_897_v, a(n_2337_v), n_897_port_4, temp_12578);
  wire [`W-1:0] temp_12579;
  spice_transistor_nmos t8862(v(clk_v), n_899_v, a(n_2335_v), n_899_port_4, temp_12579);
  spice_transistor_nmos t8863(n_1799_v, n_752_v, reg_pcl3_v, n_752_port_3, reg_pcl3_port_2);
  spice_transistor_nmos t8867(n_1800_v, reg_r3_v, n_752_v, reg_r3_port_2, n_752_port_4);
  spice_transistor_nmos t8872(n_654_v, n_753_v, reg_z3_v, n_753_port_12, reg_z3_port_2);
  spice_transistor_nmos t8875(n_657_v, reg_spl3_v, n_753_v, reg_spl3_port_2, n_753_port_13);
  spice_transistor_nmos t8876(n_658_v, n_753_v, reg_iyl3_v, n_753_port_14, reg_iyl3_port_2);
  spice_transistor_nmos t8880(n_661_v, reg_ixl3_v, n_753_v, reg_ixl3_port_2, n_753_port_15);
  spice_transistor_nmos_vdd g_8673((n_2041_v|n_795_v), n_779_v, n_779_port_8);
  spice_transistor_nmos_vdd g_8674((n_2367_v|n_2491_v), n_783_v, n_783_port_9);
  spice_transistor_nmos_vdd g_8675((n_1838_v|n_795_v), n_545_v, n_545_port_12);
  spice_transistor_nmos_vdd g_8676((n_795_v|n_2215_v), n_525_v, n_525_port_13);
  spice_transistor_nmos_vdd g_8677((n_2395_v|n_2555_v), n_808_v, n_808_port_9);
  spice_transistor_nmos_vdd g_8678((n_2444_v|n_2641_v), n_796_v, n_796_port_9);
  spice_transistor_nmos_vdd g_8679((n_2471_v|n_2231_v), n_803_v, n_803_port_9);
  spice_transistor_nmos_vdd g_8680((n_2181_v|n_2254_v), n_755_v, n_755_port_8);
  spice_transistor_nmos_vdd g_8681((n_2561_v|n_2594_v), n_836_v, n_836_port_9);
  spice_transistor_nmos_vdd g_8682((n_1751_v|v(clk_v)), n_681_v, n_681_port_6);
  spice_transistor_nmos_vdd g_8683((n_2665_v|n_2685_v), n_839_v, n_839_port_8);
  spice_transistor_nmos_vdd g_8684((n_2010_v|n_795_v), n_770_v, n_770_port_6);
  spice_transistor_nmos_vdd g_8685((n_821_v|n_822_v), n_1005_v, n_1005_port_6);
  spice_transistor_nmos_vdd g_8686((n_2321_v|n_2326_v), n_772_v, n_772_port_9);
  spice_transistor_nmos_gnd g_8688((n_135_v|n_188_v|n_95_v), n_181_v, n_181_port_7);
  spice_transistor_nmos_gnd g_8742((n_1049_v|v(n_1053_v)|n_91_v), n_75_v, n_75_port_6);
  spice_transistor_nmos_gnd g_8747((n_74_v|v(n_75_v)), n_1053_v, n_1053_port_6);
  spice_transistor_nmos_gnd g_8857((n_1141_v|v(n_128_v)), n_120_v, n_120_port_9);
  spice_transistor_nmos_gnd g_8940((n_1759_v|v(n_1783_v)), n_687_v, n_687_port_6);
  spice_transistor_nmos_gnd g_8941((v(n_687_v)|n_648_v), n_1783_v, n_1783_port_6);
  spice_transistor_nmos_gnd g_8975((v(n_1072_v)|n_131_v|n_111_v), n_86_v, n_86_port_7);
  spice_transistor_nmos_gnd g_9099((v(n_1126_v)|n_1112_v|n_135_v|n_95_v|n_188_v), n_143_v, n_143_port_7);
  spice_transistor_nmos_gnd g_9155((n_2216_v|n_2274_v), n_755_v, n_755_port_9);
  spice_transistor_nmos_gnd g_9162((n_2228_v|n_2490_v), n_803_v, n_803_port_10);
  spice_transistor_nmos_gnd g_9182((n_2297_v|n_2341_v), n_772_v, n_772_port_10);
  spice_transistor_nmos_gnd g_9192((n_131_v|v(n_1076_v)|n_111_v), n_81_v, n_81_port_7);
  spice_transistor_nmos_gnd g_9200((v(n_84_v)|n_111_v|n_131_v), n_85_v, n_85_port_8);
  spice_transistor_nmos_gnd g_9203((n_2385_v|n_2508_v), n_783_v, n_783_port_10);
  spice_transistor_nmos_gnd g_9204((n_2392_v|n_2528_v), n_808_v, n_808_port_10);
  spice_transistor_nmos_gnd g_9210((n_112_v|v(n_86_v)), n_1072_v, n_1072_port_7);
  spice_transistor_nmos_gnd g_9212((n_2417_v|n_2672_v), n_796_v, n_796_port_10);
  spice_transistor_nmos_gnd g_9218((n_1087_v|v(n_81_v)), n_1076_v, n_1076_port_7);
  spice_transistor_nmos_gnd g_9263((n_2558_v|n_2611_v), n_836_v, n_836_port_10);
  spice_transistor_nmos_gnd g_9296((n_2634_v|n_2684_v), n_839_v, n_839_port_9);
  spice_transistor_nmos_gnd g_9394((v(n_1220_v)|n_171_v), n_1204_v, n_1204_port_5);
  spice_transistor_nmos_vdd g_9433((n_608_v&v(clk_v)), n_785_v, n_785_port_17);
  spice_transistor_nmos_vdd g_9434((n_608_v&v(clk_v)), n_799_v, n_799_port_17);
  spice_transistor_nmos_vdd g_9435((n_608_v&v(clk_v)), n_914_v, n_914_port_17);
  spice_transistor_nmos_vdd g_9436((n_608_v&v(clk_v)), n_708_v, n_708_port_17);
  spice_transistor_nmos_vdd g_9437((n_608_v&v(clk_v)), n_923_v, n_923_port_17);
  spice_transistor_nmos_vdd g_9438((n_608_v&v(clk_v)), n_715_v, n_715_port_17);
  spice_transistor_nmos_vdd g_9439((n_608_v&v(clk_v)), n_807_v, n_807_port_15);
  spice_transistor_nmos_vdd g_9440((n_821_v&n_822_v), n_918_v, n_918_port_5);
  spice_transistor_nmos_vdd g_9441((n_608_v&v(clk_v)), n_934_v, n_934_port_15);
  spice_transistor_nmos_vdd g_9442((n_608_v&v(clk_v)), n_809_v, n_809_port_15);
  spice_transistor_nmos_vdd g_9443((n_608_v&v(clk_v)), n_935_v, n_935_port_15);
  spice_transistor_nmos_vdd g_9444((n_608_v&v(clk_v)), n_732_v, n_732_port_15);
  spice_transistor_nmos_vdd g_9445((n_608_v&v(clk_v)), n_949_v, n_949_port_17);
  spice_transistor_nmos_vdd g_9446((n_608_v&v(clk_v)), n_834_v, n_834_port_17);
  spice_transistor_nmos_vdd g_9447((n_608_v&v(clk_v)), n_959_v, n_959_port_17);
  spice_transistor_nmos_vdd g_9448((n_608_v&v(clk_v)), n_738_v, n_738_port_15);
  spice_transistor_nmos_vdd g_9449((n_608_v&v(clk_v)), n_847_v, n_847_port_17);
  spice_transistor_nmos_vdd g_9450((n_608_v&v(clk_v)), n_970_v, n_970_port_15);
  spice_transistor_nmos_vdd g_9451((n_608_v&v(clk_v)), n_864_v, n_864_port_15);
  spice_transistor_nmos_vdd g_9452((n_608_v&v(clk_v)), n_973_v, n_973_port_15);
  spice_transistor_nmos_vdd g_9453((n_608_v&v(clk_v)), n_745_v, n_745_port_17);
  spice_transistor_nmos_vdd g_9454((n_608_v&v(clk_v)), n_870_v, n_870_port_15);
  spice_transistor_nmos_vdd g_9455((n_608_v&v(clk_v)), n_980_v, n_980_port_17);
  spice_transistor_nmos_vdd g_9456((n_608_v&v(clk_v)), n_753_v, n_753_port_17);
  spice_transistor_nmos_vdd g_9457((n_608_v&v(clk_v)), n_985_v, n_985_port_17);
  spice_transistor_nmos_vdd g_9458((n_822_v&n_821_v), n_988_v, n_988_port_5);
  spice_transistor_nmos_vdd g_9459((n_821_v&n_822_v), n_867_v, n_867_port_5);
  spice_transistor_nmos_vdd g_9460((n_608_v&v(clk_v)), n_880_v, n_880_port_17);
  spice_transistor_nmos_vdd g_9461((n_608_v&v(clk_v)), n_999_v, n_999_port_15);
  spice_transistor_nmos_vdd g_9462((n_608_v&v(clk_v)), n_775_v, n_775_port_15);
  spice_transistor_nmos_vdd g_9463((n_608_v&v(clk_v)), n_886_v, n_886_port_17);
  spice_transistor_nmos_vdd g_9464((n_608_v&v(clk_v)), n_776_v, n_776_port_15);
  spice_transistor_nmos_vdd g_9465((n_608_v&v(clk_v)), n_902_v, n_902_port_15);
  spice_transistor_nmos_vdd g_9466((n_608_v&v(clk_v)), n_702_v, n_702_port_15);
  spice_transistor_nmos_vdd g_9467((n_608_v&v(clk_v)), n_906_v, n_906_port_15);
  spice_transistor_nmos_gnd g_9484((m6_v&n_469_v), n_1466_v, n_1466_port_4);
  spice_transistor_nmos_gnd g_9504((v(n_1466_v)&n_431_v), n_1498_v, n_1498_port_3);
  spice_transistor_nmos_gnd g_9511((n_474_v&n_1501_v), n_475_v, n_475_port_7);
  spice_transistor_nmos_gnd g_9870((v(n_359_v)&(n_1343_v|v(clk_v))), n_328_v, n_328_port_3);
  spice_transistor_nmos_gnd g_9871((v(n_1129_v)&(v(clk_v)|n_93_v)), n_132_v, n_132_port_5);
  spice_transistor_nmos_gnd g_9874((v(n_1271_v)&(v(clk_v)|n_246_v)), n_225_v, n_225_port_3);
  spice_transistor_nmos_gnd g_9880((v(n_225_v)&(n_1315_v|v(clk_v))), n_1271_v, n_1271_port_6);
  spice_transistor_nmos_gnd g_9881((v(n_1383_v)&(v(clk_v)|n_1391_v)), n_384_v, n_384_port_4);
  spice_transistor_nmos_gnd g_9886((v(n_132_v)&(n_1123_v|v(clk_v))), n_1129_v, n_1129_port_6);
  spice_transistor_nmos_gnd g_9887((v(n_223_v)&(n_1314_v|v(clk_v))), n_1184_v, n_1184_port_4);
  spice_transistor_nmos_gnd g_9888((v(n_1184_v)&(n_208_v|v(clk_v))), n_223_v, n_223_port_6);
  spice_transistor_nmos_gnd g_9890((v(n_1090_v)&(v(clk_v)|n_1106_v)), n_89_v, n_89_port_5);
  spice_transistor_nmos g_9891((n_650_v&n_1749_v), n_545_v, n_681_v, n_545_port_14, n_681_port_7);
  spice_transistor_nmos g_9892((n_650_v&n_1750_v), n_681_v, n_525_v, n_681_port_8, n_525_port_15);
  wire [`W-1:0] temp_12580;
  spice_transistor_nmos g_9894((n_650_v&n_1752_v), n_681_v, a(n_635_v), n_681_port_9, temp_12580);
  spice_transistor_nmos_gnd g_9897((v(n_89_v)&(n_1105_v|v(clk_v))), n_1090_v, n_1090_port_4);
  spice_transistor_nmos_gnd g_9898((v(n_1586_v)&(n_1563_v|v(clk_v))), n_541_v, n_541_port_3);
  spice_transistor_nmos_gnd g_9900((v(n_408_v)&(n_1404_v|v(clk_v))), n_1405_v, n_1405_port_3);
  spice_transistor_nmos_gnd g_9901((v(n_541_v)&(v(clk_v)|n_1562_v)), n_1586_v, n_1586_port_6);
  spice_transistor_nmos_gnd g_9903((v(n_244_v)&(n_1306_v|v(clk_v))), n_1327_v, n_1327_port_3);
  spice_transistor_nmos_gnd g_9907((v(n_1327_v)&(v(clk_v)|n_1307_v)), n_244_v, n_244_port_8);
  spice_transistor_nmos_gnd g_9911((v(n_127_v)&(n_1143_v|v(clk_v))), n_118_v, n_118_port_7);
  spice_transistor_nmos_gnd g_9916((v(n_94_v)&(v(clk_v)|n_1066_v)), n_1092_v, n_1092_port_5);
  spice_transistor_nmos_gnd g_9917((v(n_1098_v)&(v(clk_v)|n_1111_v)), n_92_v, n_92_port_7);
  spice_transistor_nmos_gnd g_9919((v(n_1092_v)&(n_80_v|v(clk_v))), n_94_v, n_94_port_6);
  spice_transistor_nmos_gnd g_9920((v(n_57_v)&(v(n_56_v)|v(clk_v))), n_67_v, n_67_port_5);
  spice_transistor_nmos_gnd g_9923((v(n_161_v)&(v(clk_v)|n_1190_v)), n_1170_v, n_1170_port_5);
  spice_transistor_nmos_gnd g_9927((_t2_v&(v(n_190_v)&m2_v)), n_1300_v, n_1300_port_3);
  spice_transistor_nmos_gnd g_9928((v(n_146_v)&(n_167_v|v(clk_v))), n_147_v, n_147_port_5);
  spice_transistor_nmos_gnd g_9936((v(n_1405_v)&(v(clk_v)|n_1410_v)), n_408_v, n_408_port_6);
  spice_transistor_nmos_gnd g_9943((v(n_328_v)&(v(clk_v)|n_1357_v)), n_359_v, n_359_port_6);
  spice_transistor_nmos_gnd g_9944((v(n_118_v)&(n_1153_v|v(clk_v))), n_127_v, n_127_port_6);
  spice_transistor_nmos_gnd g_9960((v(n_1051_v)&(n_1050_v|v(clk_v))), n_61_v, n_61_port_5);
  spice_transistor_nmos_gnd g_9968((v(n_176_v)&(v(n_1168_v)|v(clk_v))), n_1217_v, n_1217_port_4);
  spice_transistor_nmos_gnd g_9973((v(n_61_v)&(v(clk_v)|n_83_v)), n_1051_v, n_1051_port_6);
  spice_transistor_nmos_gnd g_9984((v(n_1649_v)&(v(clk_v)|n_577_v)), n_617_v, n_617_port_5);
  spice_transistor_nmos_gnd g_9995((v(n_617_v)&(v(clk_v)|n_685_v|n_589_v)), n_1649_v, n_1649_port_4);
  spice_transistor_nmos_gnd g_10038((v(n_62_v)&(v(clk_v)|n_1055_v)), n_1044_v, n_1044_port_3);
  spice_transistor_nmos_gnd g_10048((v(n_1170_v)&(n_1201_v|v(clk_v))), n_161_v, n_161_port_4);
  spice_transistor_nmos_gnd g_10058((v(n_67_v)&(v(clk_v)|v(n_68_v))), n_57_v, n_57_port_6);
  spice_transistor_nmos_gnd g_10059((v(n_384_v)&(v(clk_v)|n_1384_v)), n_1383_v, n_1383_port_4);
  spice_transistor_nmos_gnd g_10061((v(n_1044_v)&(v(clk_v)|n_1041_v)), n_62_v, n_62_port_6);
  spice_transistor_nmos_gnd g_10068((v(n_147_v)&(n_1177_v|v(clk_v))), n_146_v, n_146_port_4);
  spice_transistor_nmos_gnd g_10077((v(n_92_v)&(n_129_v|v(clk_v))), n_1098_v, n_1098_port_4);
  spice_transistor_nmos_gnd g_10115((v(n_175_v)|(n_1152_v&n_162_v)), n_1225_v, n_1225_port_7);
  spice_transistor_nmos_gnd g_10116((v(n_1218_v)|(n_1238_v&n_162_v)), n_1228_v, n_1228_port_7);
  spice_transistor_nmos_gnd g_10120((v(n_77_v)|(v(n_1051_v)&v(clk_v))), n_1060_v, n_1060_port_5);
  spice_transistor_nmos_gnd g_10128((v(n_197_v)|(v(n_136_v)&n_1265_v)), n_185_v, n_185_port_7);
  spice_transistor_nmos_gnd g_10130((v(n_1060_v)|(v(n_61_v)&v(clk_v))), n_77_v, n_77_port_8);
  spice_transistor_nmos_gnd g_10131((n_220_v|(n_232_v&n_1256_v)), n_1232_v, n_1232_port_5);
  spice_transistor_nmos_gnd g_10133((v(n_185_v)|(v(n_139_v)&n_1265_v)), n_197_v, n_197_port_6);
  spice_transistor_nmos_gnd g_10134((v(n_56_v)|(v(n_58_v)&n_59_v)), n_68_v, n_68_port_9);
  spice_transistor_nmos_gnd g_10135((v(n_1095_v)|(v(n_1092_v)&v(clk_v))), n_1079_v, n_1079_port_5);
  spice_transistor_nmos_gnd g_10139((v(n_70_v)|(v(n_67_v)&v(clk_v))), n_73_v, n_73_port_6);
  spice_transistor_nmos_gnd g_10140((v(n_73_v)|(v(n_57_v)&v(clk_v))), n_70_v, n_70_port_7);
  spice_transistor_nmos_gnd g_10143((v(n_216_v)|(v(clk_v)&(_t1_v&m1_v))), n_1320_v, n_1320_port_5);
  spice_transistor_nmos_gnd g_10144((v(n_240_v)|(n_211_v&v(clk_v))), n_214_v, n_214_port_5);
  spice_transistor_nmos_gnd g_10146((v(n_214_v)|(n_1333_v&v(clk_v))), n_240_v, n_240_port_8);
  spice_transistor_nmos_gnd g_10151((v(n_1313_v)|(v(n_1302_v)&v(clk_v))), n_241_v, n_241_port_7);
  spice_transistor_nmos_gnd g_10154((v(n_1320_v)|(v(clk_v)&(n_66_v|_t3_v))), n_216_v, n_216_port_8);
  spice_transistor_nmos_gnd g_10155((v(n_241_v)|(v(clk_v)&(m4_v|m1_v))), n_1313_v, n_1313_port_6);
  spice_transistor_nmos_gnd g_10157((v(n_1701_v)|(n_1731_v&n_1722_v)), ex_dehl0_v, ex_dehl0_port_9);
  spice_transistor_nmos_gnd g_10158((v(n_1702_v)|(n_1728_v&n_1719_v)), ex_dehl1_v, ex_dehl1_port_9);
  spice_transistor_nmos_gnd g_10159((v(ex_dehl1_v)|(n_1727_v&n_1719_v)), n_1702_v, n_1702_port_8);
  spice_transistor_nmos_gnd g_10160((v(ex_dehl0_v)|(n_1730_v&n_1722_v)), n_1701_v, n_1701_port_8);
  spice_transistor_nmos_gnd g_10162((n_55_v|(n_59_v&v(n_1043_v))), n_58_v, n_58_port_8);
  spice_transistor_nmos_gnd g_10164((v(n_1161_v)|(v(clk_v)&(n_141_v&n_54_v))), n_1168_v, n_1168_port_8);
  spice_transistor_nmos_gnd g_10166((v(ex_af_v)|(n_1768_v&n_639_v)), n_633_v, n_633_port_9);
  spice_transistor_nmos_gnd g_10167((v(n_633_v)|(n_1767_v&n_639_v)), ex_af_v, ex_af_port_10);
  spice_transistor_nmos_gnd g_10168((v(n_124_v)|(n_145_v&v(clk_v))), n_1080_v, n_1080_port_8);
  spice_transistor_nmos_gnd g_10169((v(n_1773_v)|(n_1771_v&n_1716_v)), ex_bcdehl_v, ex_bcdehl_port_8);
  spice_transistor_nmos_gnd g_10170((v(ex_bcdehl_v)|(n_1772_v&n_1716_v)), n_1773_v, n_1773_port_9);
  spice_transistor_nmos_gnd g_10171((v(n_1168_v)|(n_1165_v&v(clk_v))), n_1161_v, n_1161_port_9);
  spice_transistor_nmos_gnd g_10172((v(n_259_v)|(n_1334_v&n_162_v)), n_1341_v, n_1341_port_5);
  spice_transistor_nmos_gnd g_10174((v(n_139_v)|(v(n_1129_v)&v(clk_v))), n_136_v, n_136_port_10);
  spice_transistor_nmos_gnd g_10176((v(n_1341_v)|(n_126_v&n_162_v)), n_259_v, n_259_port_8);
  spice_transistor_nmos_gnd g_10178((v(n_143_v)|(n_97_v&n_122_v)), n_1126_v, n_1126_port_8);
  spice_transistor_nmos_gnd g_10179((v(n_150_v)|(n_114_v&n_122_v)), n_149_v, n_149_port_8);
  spice_transistor_nmos_gnd g_10181((v(n_1079_v)|(v(n_94_v)&v(clk_v))), n_1095_v, n_1095_port_8);
  spice_transistor_nmos_gnd g_10182((v(n_148_v)|(n_106_v&n_122_v)), n_1171_v, n_1171_port_7);
  spice_transistor_nmos_gnd g_10184((v(n_1178_v)|(n_1137_v&n_162_v)), n_140_v, n_140_port_7);
  spice_transistor_nmos_gnd g_10187((v(n_140_v)|(n_1144_v&n_162_v)), n_1178_v, n_1178_port_6);
  spice_transistor_nmos_gnd g_10189((v(n_136_v)|(v(n_132_v)&v(clk_v))), n_139_v, n_139_port_12);
  spice_transistor_nmos_gnd g_10192((v(n_98_v)|(v(clk_v)&(n_125_v&_t3_v))), n_1077_v, n_1077_port_8);
  spice_transistor_nmos_gnd g_10196((v(n_172_v)|(v(n_136_v)&n_153_v)), n_157_v, n_157_port_8);
  spice_transistor_nmos_gnd g_10199((v(n_169_v)|(n_1151_v&n_162_v)), n_1221_v, n_1221_port_7);
  spice_transistor_nmos_gnd g_10200((v(n_1221_v)|(n_158_v&n_162_v)), n_169_v, n_169_port_6);
  spice_transistor_nmos_gnd g_10201((n_65_v|(v(n_1217_v)&(v(clk_v)|v(n_1161_v)))), n_176_v, n_176_port_10);
  spice_transistor_nmos_gnd g_10203((v(n_1225_v)|(n_1179_v&n_162_v)), n_175_v, n_175_port_6);
  spice_transistor_nmos_gnd g_10204((v(n_1228_v)|(n_1213_v&n_162_v)), n_1218_v, n_1218_port_6);
  spice_transistor_nmos_gnd g_10213(((n_1234_v|v(n_1204_v))|(_t1_v&v(clk_v))), n_1220_v, n_1220_port_10);
  spice_transistor_nmos_gnd g_10214(((n_95_v|v(n_157_v))|(n_153_v&(n_174_v&v(n_139_v)))), n_172_v, n_172_port_8);
  spice_transistor_nmos_gnd g_10219(((n_55_v|v(n_68_v))|(v(n_1043_v)&n_59_v)), n_56_v, n_56_port_11);
  spice_transistor_nmos_gnd g_10220(((v(n_1080_v)|n_1081_v)|(n_1082_v&v(clk_v))), n_124_v, n_124_port_9);
  spice_transistor_nmos_gnd g_10223(((n_1128_v|v(n_120_v))|(n_1121_v&v(clk_v))), n_128_v, n_128_port_10);
  spice_transistor_nmos_gnd g_10226(((v(n_149_v)|n_95_v)|(n_1110_v&n_122_v)), n_150_v, n_150_port_11);
  spice_transistor_nmos_gnd g_10227(((v(n_1171_v)|n_95_v)|(n_1127_v&n_122_v)), n_148_v, n_148_port_13);
  spice_transistor_nmos_gnd g_10229(((n_1083_v|v(n_85_v))|(n_1084_v&v(clk_v))), n_84_v, n_84_port_10);
  spice_transistor_nmos_gnd g_10230(((n_95_v|v(n_1077_v))|(v(clk_v)&(_t2_v|n_107_v))), n_98_v, n_98_port_8);
  spice_transistor_nmos_vdd g_10313((v(n_562_v)&(n_1632_v|(v(n_562_v)&(n_66_v&v(clk_v))))), vss_v, vss_port_5680);

  spice_pullup pullup_6578(n_61_v, n_61_port_3);
  spice_pullup pullup_6579(n_62_v, n_62_port_3);
  spice_pullup pullup_6582(n_75_v, n_75_port_5);
  spice_pullup pullup_6584(n_77_v, n_77_port_5);
  spice_pullup pullup_6585(n_81_v, n_81_port_6);
  spice_pullup pullup_6586(n_89_v, n_89_port_4);
  spice_pullup pullup_6588(n_92_v, n_92_port_4);
  spice_pullup pullup_6591(n_118_v, n_118_port_4);
  spice_pullup pullup_6592(n_120_v, n_120_port_5);
  spice_pullup pullup_6593(n_127_v, n_127_port_3);
  spice_pullup pullup_6594(n_128_v, n_128_port_6);
  spice_pullup pullup_6595(n_132_v, n_132_port_3);
  spice_pullup pullup_6596(n_136_v, n_136_port_5);
  spice_pullup pullup_6597(n_139_v, n_139_port_5);
  spice_pullup pullup_6598(n_140_v, n_140_port_5);
  spice_pullup pullup_6600(n_146_v, n_146_port_2);
  spice_pullup pullup_6601(n_147_v, n_147_port_4);
  spice_pullup pullup_6605(n_157_v, n_157_port_4);
  spice_pullup pullup_6607(n_161_v, n_161_port_2);
  spice_pullup pullup_6609(n_169_v, n_169_port_3);
  spice_pullup pullup_6610(n_172_v, n_172_port_4);
  spice_pullup pullup_6612(n_175_v, n_175_port_3);
  spice_pullup pullup_6613(n_176_v, n_176_port_5);
  spice_pullup pullup_6615(n_185_v, n_185_port_5);
  spice_pullup pullup_6617(n_190_v, n_190_port_3);
  spice_pullup pullup_6619(n_197_v, n_197_port_3);
  spice_pullup pullup_6627(n_214_v, n_214_port_3);
  spice_pullup pullup_6629(n_216_v, n_216_port_5);
  spice_pullup pullup_6632(n_223_v, n_223_port_3);
  spice_pullup pullup_6634(n_225_v, n_225_port_2);
  spice_pullup pullup_6640(n_240_v, n_240_port_5);
  spice_pullup pullup_6641(n_241_v, n_241_port_5);
  spice_pullup pullup_6650(n_259_v, n_259_port_5);
  spice_pullup pullup_6672(n_328_v, n_328_port_2);
  spice_pullup pullup_6687(n_56_v, n_56_port_5);
  spice_pullup pullup_6688(n_57_v, n_57_port_3);
  spice_pullup pullup_6689(n_58_v, n_58_port_4);
  spice_pullup pullup_6691(n_67_v, n_67_port_3);
  spice_pullup pullup_6692(n_68_v, n_68_port_4);
  spice_pullup pullup_6693(n_70_v, n_70_port_4);
  spice_pullup pullup_6694(n_73_v, n_73_port_4);
  spice_pullup pullup_6696(n_84_v, n_84_port_6);
  spice_pullup pullup_6697(n_85_v, n_85_port_6);
  spice_pullup pullup_6698(n_86_v, n_86_port_6);
  spice_pullup pullup_6699(n_94_v, n_94_port_3);
  spice_pullup pullup_6701(n_98_v, n_98_port_4);
  spice_pullup pullup_6709(n_124_v, n_124_port_5);
  spice_pullup pullup_6713(n_143_v, n_143_port_6);
  spice_pullup pullup_6715(n_148_v, n_148_port_6);
  spice_pullup pullup_6716(n_149_v, n_149_port_5);
  spice_pullup pullup_6717(n_150_v, n_150_port_5);
  spice_pullup pullup_6741(n_244_v, n_244_port_4);
  spice_pullup pullup_6803(n_359_v, n_359_port_3);
  spice_pullup pullup_6812(n_384_v, n_384_port_3);
  spice_pullup pullup_6824(n_408_v, n_408_port_4);
  spice_pullup pullup_6956(n_617_v, n_617_port_3);
  spice_pullup pullup_6957(ex_dehl0_v, ex_dehl0_port_5);
  spice_pullup pullup_6960(ex_dehl1_v, ex_dehl1_port_5);
  spice_pullup pullup_6963(n_633_v, n_633_port_5);
  spice_pullup pullup_6983(n_707_v, n_707_port_3);
  spice_pullup pullup_6984(n_709_v, n_709_port_5);
  spice_pullup pullup_6987(n_721_v, n_721_port_4);
  spice_pullup pullup_6988(n_722_v, n_722_port_3);
  spice_pullup pullup_6993(n_744_v, n_744_port_3);
  spice_pullup pullup_6994(n_746_v, n_746_port_5);
  spice_pullup pullup_6997(n_763_v, n_763_port_4);
  spice_pullup pullup_6998(n_769_v, n_769_port_3);
  spice_pullup pullup_7004(n_784_v, n_784_port_3);
  spice_pullup pullup_7005(n_787_v, n_787_port_5);
  spice_pullup pullup_7008(n_802_v, n_802_port_4);
  spice_pullup pullup_7009(n_804_v, n_804_port_3);
  spice_pullup pullup_7014(n_833_v, n_833_port_3);
  spice_pullup pullup_7015(n_835_v, n_835_port_3);
  spice_pullup pullup_7019(n_856_v, n_856_port_5);
  spice_pullup pullup_7020(n_857_v, n_857_port_3);
  spice_pullup pullup_7037(n_541_v, n_541_port_2);
  spice_pullup pullup_7059(ex_af_v, ex_af_port_5);
  spice_pullup pullup_7075(n_687_v, n_687_port_5);
  spice_pullup pullup_7079(n_700_v, n_700_port_3);
  spice_pullup pullup_7088(n_728_v, n_728_port_4);
  spice_pullup pullup_7092(n_754_v, n_754_port_5);
  spice_pullup pullup_7120(n_879_v, n_879_port_3);
  spice_pullup pullup_7121(n_881_v, n_881_port_4);
  spice_pullup pullup_7126(n_892_v, n_892_port_5);
  spice_pullup pullup_7127(n_893_v, n_893_port_3);
  spice_pullup pullup_7132(n_913_v, n_913_port_3);
  spice_pullup pullup_7133(n_915_v, n_915_port_4);
  spice_pullup pullup_7135(n_928_v, n_928_port_3);
  spice_pullup pullup_7136(n_929_v, n_929_port_3);
  spice_pullup pullup_7142(n_948_v, n_948_port_3);
  spice_pullup pullup_7143(n_950_v, n_950_port_5);
  spice_pullup pullup_7146(n_963_v, n_963_port_4);
  spice_pullup pullup_7147(n_964_v, n_964_port_3);
  spice_pullup pullup_7152(n_979_v, n_979_port_3);
  spice_pullup pullup_7153(n_981_v, n_981_port_3);
  spice_pullup pullup_7155(n_994_v, n_994_port_3);
  spice_pullup pullup_7163(n_861_v, n_861_port_3);
  spice_pullup pullup_7173(n_908_v, n_908_port_3);
  spice_pullup pullup_7181(n_956_v, n_956_port_4);
  spice_pullup pullup_7189(n_1001_v, n_1001_port_4);
  spice_pullup pullup_7202(n_1051_v, n_1051_port_3);
  spice_pullup pullup_7203(n_1044_v, n_1044_port_2);
  spice_pullup pullup_7206(n_1053_v, n_1053_port_4);
  spice_pullup pullup_7207(n_1060_v, n_1060_port_3);
  spice_pullup pullup_7215(n_1090_v, n_1090_port_2);
  spice_pullup pullup_7221(n_1098_v, n_1098_port_2);
  spice_pullup pullup_7227(n_1129_v, n_1129_port_3);
  spice_pullup pullup_7241(n_1168_v, n_1168_port_4);
  spice_pullup pullup_7242(n_1161_v, n_1161_port_4);
  spice_pullup pullup_7249(n_1170_v, n_1170_port_4);
  spice_pullup pullup_7251(n_1178_v, n_1178_port_3);
  spice_pullup pullup_7264(n_1218_v, n_1218_port_3);
  spice_pullup pullup_7265(n_1217_v, n_1217_port_2);
  spice_pullup pullup_7267(n_1221_v, n_1221_port_5);
  spice_pullup pullup_7268(n_1225_v, n_1225_port_5);
  spice_pullup pullup_7269(n_1228_v, n_1228_port_5);
  spice_pullup pullup_7282(n_1232_v, n_1232_port_3);
  spice_pullup pullup_7287(n_1300_v, n_1300_port_2);
  spice_pullup pullup_7292(n_1302_v, n_1302_port_2);
  spice_pullup pullup_7293(n_1320_v, n_1320_port_3);
  spice_pullup pullup_7296(n_1271_v, n_1271_port_4);
  spice_pullup pullup_7297(n_1313_v, n_1313_port_3);
  spice_pullup pullup_7298(n_1184_v, n_1184_port_3);
  spice_pullup pullup_7304(n_1332_v, n_1332_port_2);
  spice_pullup pullup_7310(n_1341_v, n_1341_port_3);
  spice_pullup pullup_7322(n_1383_v, n_1383_port_2);
  spice_pullup pullup_7335(n_1405_v, n_1405_port_2);
  spice_pullup pullup_7434(n_1649_v, n_1649_port_2);
  spice_pullup pullup_7450(n_1701_v, n_1701_port_4);
  spice_pullup pullup_7451(n_1702_v, n_1702_port_4);
  spice_pullup pullup_7468(ex_bcdehl_v, ex_bcdehl_port_5);
  spice_pullup pullup_7469(n_1773_v, n_1773_port_5);
  spice_pullup pullup_7480(n_1814_v, n_1814_port_3);
  spice_pullup pullup_7481(n_1815_v, n_1815_port_3);
  spice_pullup pullup_7482(n_1816_v, n_1816_port_3);
  spice_pullup pullup_7483(n_1817_v, n_1817_port_3);
  spice_pullup pullup_7484(n_1818_v, n_1818_port_3);
  spice_pullup pullup_7485(n_1819_v, n_1819_port_3);
  spice_pullup pullup_7486(n_1820_v, n_1820_port_3);
  spice_pullup pullup_7487(n_1821_v, n_1821_port_3);
  spice_pullup pullup_7488(n_1822_v, n_1822_port_3);
  spice_pullup pullup_7489(n_1823_v, n_1823_port_3);
  spice_pullup pullup_7490(n_1824_v, n_1824_port_3);
  spice_pullup pullup_7491(n_1825_v, n_1825_port_3);
  spice_pullup pullup_7492(n_1826_v, n_1826_port_3);
  spice_pullup pullup_7493(n_1827_v, n_1827_port_3);
  spice_pullup pullup_7500(reg_pcl0_v, reg_pcl0_port_3);
  spice_pullup pullup_7501(reg_r0_v, reg_r0_port_3);
  spice_pullup pullup_7502(reg_z0_v, reg_z0_port_3);
  spice_pullup pullup_7503(reg_spl0_v, reg_spl0_port_3);
  spice_pullup pullup_7504(reg_iyl0_v, reg_iyl0_port_3);
  spice_pullup pullup_7505(reg_ixl0_v, reg_ixl0_port_3);
  spice_pullup pullup_7506(reg_e0_v, reg_e0_port_3);
  spice_pullup pullup_7507(reg_ee0_v, reg_ee0_port_3);
  spice_pullup pullup_7508(reg_l0_v, reg_l0_port_3);
  spice_pullup pullup_7509(reg_ll0_v, reg_ll0_port_3);
  spice_pullup pullup_7510(reg_c0_v, reg_c0_port_3);
  spice_pullup pullup_7511(reg_cc0_v, reg_cc0_port_3);
  spice_pullup pullup_7512(reg_ff0_v, reg_ff0_port_3);
  spice_pullup pullup_7513(reg_f0_v, reg_f0_port_3);
  spice_pullup pullup_7519(reg_pcl1_v, reg_pcl1_port_3);
  spice_pullup pullup_7520(reg_r1_v, reg_r1_port_3);
  spice_pullup pullup_7523(reg_z1_v, reg_z1_port_3);
  spice_pullup pullup_7524(reg_spl1_v, reg_spl1_port_3);
  spice_pullup pullup_7525(reg_iyl1_v, reg_iyl1_port_3);
  spice_pullup pullup_7526(reg_ixl1_v, reg_ixl1_port_3);
  spice_pullup pullup_7527(reg_e1_v, reg_e1_port_3);
  spice_pullup pullup_7528(reg_ee1_v, reg_ee1_port_3);
  spice_pullup pullup_7529(reg_l1_v, reg_l1_port_3);
  spice_pullup pullup_7530(reg_ll1_v, reg_ll1_port_3);
  spice_pullup pullup_7531(reg_c1_v, reg_c1_port_3);
  spice_pullup pullup_7532(reg_cc1_v, reg_cc1_port_3);
  spice_pullup pullup_7533(reg_ff1_v, reg_ff1_port_3);
  spice_pullup pullup_7534(reg_f1_v, reg_f1_port_3);
  spice_pullup pullup_7536(n_1890_v, n_1890_port_3);
  spice_pullup pullup_7537(n_1891_v, n_1891_port_3);
  spice_pullup pullup_7538(n_1892_v, n_1892_port_3);
  spice_pullup pullup_7539(n_1893_v, n_1893_port_3);
  spice_pullup pullup_7540(n_1894_v, n_1894_port_3);
  spice_pullup pullup_7541(n_1895_v, n_1895_port_3);
  spice_pullup pullup_7542(n_1896_v, n_1896_port_3);
  spice_pullup pullup_7543(n_1897_v, n_1897_port_3);
  spice_pullup pullup_7544(n_1898_v, n_1898_port_3);
  spice_pullup pullup_7545(n_1899_v, n_1899_port_3);
  spice_pullup pullup_7546(n_1900_v, n_1900_port_3);
  spice_pullup pullup_7547(n_1901_v, n_1901_port_3);
  spice_pullup pullup_7548(n_1902_v, n_1902_port_3);
  spice_pullup pullup_7549(n_1903_v, n_1903_port_3);
  spice_pullup pullup_7556(n_1915_v, n_1915_port_3);
  spice_pullup pullup_7557(n_1916_v, n_1916_port_3);
  spice_pullup pullup_7558(n_1917_v, n_1917_port_3);
  spice_pullup pullup_7559(n_1918_v, n_1918_port_3);
  spice_pullup pullup_7560(n_1919_v, n_1919_port_3);
  spice_pullup pullup_7561(n_1920_v, n_1920_port_3);
  spice_pullup pullup_7562(n_1921_v, n_1921_port_3);
  spice_pullup pullup_7563(n_1922_v, n_1922_port_3);
  spice_pullup pullup_7564(n_1923_v, n_1923_port_3);
  spice_pullup pullup_7565(n_1924_v, n_1924_port_3);
  spice_pullup pullup_7566(n_1925_v, n_1925_port_3);
  spice_pullup pullup_7567(n_1926_v, n_1926_port_3);
  spice_pullup pullup_7568(n_1927_v, n_1927_port_3);
  spice_pullup pullup_7569(n_1928_v, n_1928_port_3);
  spice_pullup pullup_7576(reg_pcl2_v, reg_pcl2_port_3);
  spice_pullup pullup_7577(reg_r2_v, reg_r2_port_3);
  spice_pullup pullup_7578(reg_z2_v, reg_z2_port_3);
  spice_pullup pullup_7579(reg_spl2_v, reg_spl2_port_3);
  spice_pullup pullup_7580(reg_iyl2_v, reg_iyl2_port_3);
  spice_pullup pullup_7581(reg_ixl2_v, reg_ixl2_port_3);
  spice_pullup pullup_7582(reg_e2_v, reg_e2_port_3);
  spice_pullup pullup_7583(reg_ee2_v, reg_ee2_port_3);
  spice_pullup pullup_7584(reg_l2_v, reg_l2_port_3);
  spice_pullup pullup_7585(reg_ll2_v, reg_ll2_port_3);
  spice_pullup pullup_7586(reg_c2_v, reg_c2_port_3);
  spice_pullup pullup_7587(reg_cc2_v, reg_cc2_port_3);
  spice_pullup pullup_7588(reg_ff2_v, reg_ff2_port_3);
  spice_pullup pullup_7589(reg_f2_v, reg_f2_port_3);
  spice_pullup pullup_7594(reg_pcl3_v, reg_pcl3_port_3);
  spice_pullup pullup_7595(reg_r3_v, reg_r3_port_3);
  spice_pullup pullup_7597(reg_z3_v, reg_z3_port_3);
  spice_pullup pullup_7598(reg_spl3_v, reg_spl3_port_3);
  spice_pullup pullup_7599(reg_iyl3_v, reg_iyl3_port_3);
  spice_pullup pullup_7600(reg_ixl3_v, reg_ixl3_port_3);
  spice_pullup pullup_7601(reg_e3_v, reg_e3_port_3);
  spice_pullup pullup_7602(reg_ee3_v, reg_ee3_port_3);
  spice_pullup pullup_7603(reg_l3_v, reg_l3_port_3);
  spice_pullup pullup_7604(reg_ll3_v, reg_ll3_port_3);
  spice_pullup pullup_7605(reg_c3_v, reg_c3_port_3);
  spice_pullup pullup_7606(reg_cc3_v, reg_cc3_port_3);
  spice_pullup pullup_7607(reg_ff3_v, reg_ff3_port_3);
  spice_pullup pullup_7608(reg_f3_v, reg_f3_port_3);
  spice_pullup pullup_7612(n_1996_v, n_1996_port_3);
  spice_pullup pullup_7613(n_1997_v, n_1997_port_3);
  spice_pullup pullup_7614(n_1998_v, n_1998_port_3);
  spice_pullup pullup_7615(n_1999_v, n_1999_port_3);
  spice_pullup pullup_7616(n_2000_v, n_2000_port_3);
  spice_pullup pullup_7617(n_2001_v, n_2001_port_3);
  spice_pullup pullup_7618(n_2002_v, n_2002_port_3);
  spice_pullup pullup_7619(n_2003_v, n_2003_port_3);
  spice_pullup pullup_7620(n_2004_v, n_2004_port_3);
  spice_pullup pullup_7621(n_2005_v, n_2005_port_3);
  spice_pullup pullup_7622(n_2006_v, n_2006_port_3);
  spice_pullup pullup_7623(n_2007_v, n_2007_port_3);
  spice_pullup pullup_7624(n_2008_v, n_2008_port_3);
  spice_pullup pullup_7625(n_2009_v, n_2009_port_3);
  spice_pullup pullup_7632(n_2019_v, n_2019_port_3);
  spice_pullup pullup_7633(n_2020_v, n_2020_port_3);
  spice_pullup pullup_7634(n_2021_v, n_2021_port_3);
  spice_pullup pullup_7635(n_2022_v, n_2022_port_3);
  spice_pullup pullup_7636(n_2023_v, n_2023_port_3);
  spice_pullup pullup_7637(n_2024_v, n_2024_port_3);
  spice_pullup pullup_7638(n_2025_v, n_2025_port_3);
  spice_pullup pullup_7639(n_2026_v, n_2026_port_3);
  spice_pullup pullup_7640(n_2027_v, n_2027_port_3);
  spice_pullup pullup_7641(n_2028_v, n_2028_port_3);
  spice_pullup pullup_7642(n_2029_v, n_2029_port_3);
  spice_pullup pullup_7643(n_2030_v, n_2030_port_3);
  spice_pullup pullup_7644(n_2031_v, n_2031_port_3);
  spice_pullup pullup_7645(n_2032_v, n_2032_port_3);
  spice_pullup pullup_7651(reg_pcl4_v, reg_pcl4_port_3);
  spice_pullup pullup_7652(reg_r4_v, reg_r4_port_3);
  spice_pullup pullup_7653(reg_z4_v, reg_z4_port_3);
  spice_pullup pullup_7654(reg_spl4_v, reg_spl4_port_3);
  spice_pullup pullup_7655(reg_iyl4_v, reg_iyl4_port_3);
  spice_pullup pullup_7656(reg_ixl4_v, reg_ixl4_port_3);
  spice_pullup pullup_7657(reg_e4_v, reg_e4_port_3);
  spice_pullup pullup_7658(reg_ee4_v, reg_ee4_port_3);
  spice_pullup pullup_7659(reg_l4_v, reg_l4_port_3);
  spice_pullup pullup_7660(reg_ll4_v, reg_ll4_port_3);
  spice_pullup pullup_7661(reg_c4_v, reg_c4_port_3);
  spice_pullup pullup_7662(reg_cc4_v, reg_cc4_port_3);
  spice_pullup pullup_7663(reg_ff4_v, reg_ff4_port_3);
  spice_pullup pullup_7664(reg_f4_v, reg_f4_port_3);
  spice_pullup pullup_7669(reg_pcl5_v, reg_pcl5_port_3);
  spice_pullup pullup_7670(reg_r5_v, reg_r5_port_3);
  spice_pullup pullup_7672(reg_z5_v, reg_z5_port_3);
  spice_pullup pullup_7673(reg_spl5_v, reg_spl5_port_3);
  spice_pullup pullup_7674(reg_iyl5_v, reg_iyl5_port_3);
  spice_pullup pullup_7675(reg_ixl5_v, reg_ixl5_port_3);
  spice_pullup pullup_7676(reg_e5_v, reg_e5_port_3);
  spice_pullup pullup_7677(reg_ee5_v, reg_ee5_port_3);
  spice_pullup pullup_7678(reg_l5_v, reg_l5_port_3);
  spice_pullup pullup_7679(reg_ll5_v, reg_ll5_port_3);
  spice_pullup pullup_7680(reg_c5_v, reg_c5_port_3);
  spice_pullup pullup_7681(reg_cc5_v, reg_cc5_port_3);
  spice_pullup pullup_7682(reg_ff5_v, reg_ff5_port_3);
  spice_pullup pullup_7683(reg_f5_v, reg_f5_port_3);
  spice_pullup pullup_7686(n_2094_v, n_2094_port_3);
  spice_pullup pullup_7687(n_2095_v, n_2095_port_3);
  spice_pullup pullup_7688(n_2096_v, n_2096_port_3);
  spice_pullup pullup_7689(n_2097_v, n_2097_port_3);
  spice_pullup pullup_7690(n_2098_v, n_2098_port_3);
  spice_pullup pullup_7691(n_2099_v, n_2099_port_3);
  spice_pullup pullup_7692(n_2100_v, n_2100_port_3);
  spice_pullup pullup_7693(n_2101_v, n_2101_port_3);
  spice_pullup pullup_7694(n_2102_v, n_2102_port_3);
  spice_pullup pullup_7695(n_2103_v, n_2103_port_3);
  spice_pullup pullup_7696(n_2104_v, n_2104_port_3);
  spice_pullup pullup_7697(n_2105_v, n_2105_port_3);
  spice_pullup pullup_7698(n_2106_v, n_2106_port_3);
  spice_pullup pullup_7699(n_2107_v, n_2107_port_3);
  spice_pullup pullup_7705(n_2119_v, n_2119_port_3);
  spice_pullup pullup_7706(n_2120_v, n_2120_port_3);
  spice_pullup pullup_7707(n_2121_v, n_2121_port_3);
  spice_pullup pullup_7708(n_2122_v, n_2122_port_3);
  spice_pullup pullup_7709(n_2123_v, n_2123_port_3);
  spice_pullup pullup_7710(n_2124_v, n_2124_port_3);
  spice_pullup pullup_7711(n_2125_v, n_2125_port_3);
  spice_pullup pullup_7712(n_2126_v, n_2126_port_3);
  spice_pullup pullup_7713(n_2127_v, n_2127_port_3);
  spice_pullup pullup_7714(n_2128_v, n_2128_port_3);
  spice_pullup pullup_7715(n_2129_v, n_2129_port_3);
  spice_pullup pullup_7716(n_2130_v, n_2130_port_3);
  spice_pullup pullup_7717(n_2131_v, n_2131_port_3);
  spice_pullup pullup_7718(n_2132_v, n_2132_port_3);
  spice_pullup pullup_7725(reg_pcl6_v, reg_pcl6_port_3);
  spice_pullup pullup_7726(reg_r6_v, reg_r6_port_3);
  spice_pullup pullup_7727(reg_z6_v, reg_z6_port_3);
  spice_pullup pullup_7728(reg_spl6_v, reg_spl6_port_3);
  spice_pullup pullup_7729(reg_iyl6_v, reg_iyl6_port_3);
  spice_pullup pullup_7730(reg_ixl6_v, reg_ixl6_port_3);
  spice_pullup pullup_7731(reg_e6_v, reg_e6_port_3);
  spice_pullup pullup_7732(reg_ee6_v, reg_ee6_port_3);
  spice_pullup pullup_7733(reg_l6_v, reg_l6_port_3);
  spice_pullup pullup_7734(reg_ll6_v, reg_ll6_port_3);
  spice_pullup pullup_7735(reg_c6_v, reg_c6_port_3);
  spice_pullup pullup_7736(reg_cc6_v, reg_cc6_port_3);
  spice_pullup pullup_7737(reg_ff6_v, reg_ff6_port_3);
  spice_pullup pullup_7738(reg_f6_v, reg_f6_port_3);
  spice_pullup pullup_7742(reg_pcl7_v, reg_pcl7_port_3);
  spice_pullup pullup_7743(reg_r7_v, reg_r7_port_3);
  spice_pullup pullup_7745(reg_z7_v, reg_z7_port_3);
  spice_pullup pullup_7746(reg_spl7_v, reg_spl7_port_3);
  spice_pullup pullup_7747(reg_iyl7_v, reg_iyl7_port_3);
  spice_pullup pullup_7748(reg_ixl7_v, reg_ixl7_port_3);
  spice_pullup pullup_7749(reg_e7_v, reg_e7_port_3);
  spice_pullup pullup_7750(reg_ee7_v, reg_ee7_port_3);
  spice_pullup pullup_7751(reg_l7_v, reg_l7_port_3);
  spice_pullup pullup_7752(reg_ll7_v, reg_ll7_port_3);
  spice_pullup pullup_7753(reg_c7_v, reg_c7_port_3);
  spice_pullup pullup_7754(reg_cc7_v, reg_cc7_port_3);
  spice_pullup pullup_7755(reg_ff7_v, reg_ff7_port_3);
  spice_pullup pullup_7756(reg_f7_v, reg_f7_port_3);
  spice_pullup pullup_7759(n_2196_v, n_2196_port_3);
  spice_pullup pullup_7760(n_2197_v, n_2197_port_3);
  spice_pullup pullup_7761(n_2198_v, n_2198_port_3);
  spice_pullup pullup_7762(n_2199_v, n_2199_port_3);
  spice_pullup pullup_7763(n_2200_v, n_2200_port_3);
  spice_pullup pullup_7764(n_2201_v, n_2201_port_3);
  spice_pullup pullup_7765(n_2202_v, n_2202_port_3);
  spice_pullup pullup_7766(n_2203_v, n_2203_port_3);
  spice_pullup pullup_7767(n_2204_v, n_2204_port_3);
  spice_pullup pullup_7768(n_2205_v, n_2205_port_3);
  spice_pullup pullup_7769(n_2206_v, n_2206_port_3);
  spice_pullup pullup_7770(n_2207_v, n_2207_port_3);
  spice_pullup pullup_7771(n_2208_v, n_2208_port_3);
  spice_pullup pullup_7772(n_2209_v, n_2209_port_3);
  spice_pullup pullup_7779(n_2232_v, n_2232_port_3);
  spice_pullup pullup_7780(n_2233_v, n_2233_port_3);
  spice_pullup pullup_7781(n_2234_v, n_2234_port_3);
  spice_pullup pullup_7782(n_2235_v, n_2235_port_3);
  spice_pullup pullup_7783(n_2236_v, n_2236_port_3);
  spice_pullup pullup_7784(n_2237_v, n_2237_port_3);
  spice_pullup pullup_7785(n_2238_v, n_2238_port_3);
  spice_pullup pullup_7786(n_2239_v, n_2239_port_3);
  spice_pullup pullup_7787(n_2240_v, n_2240_port_3);
  spice_pullup pullup_7788(n_2241_v, n_2241_port_3);
  spice_pullup pullup_7789(n_2242_v, n_2242_port_3);
  spice_pullup pullup_7790(n_2243_v, n_2243_port_3);
  spice_pullup pullup_7791(n_2244_v, n_2244_port_3);
  spice_pullup pullup_7792(n_2245_v, n_2245_port_3);
  spice_pullup pullup_7798(reg_pch0_v, reg_pch0_port_3);
  spice_pullup pullup_7799(reg_i0_v, reg_i0_port_3);
  spice_pullup pullup_7800(reg_w0_v, reg_w0_port_3);
  spice_pullup pullup_7801(reg_sph0_v, reg_sph0_port_3);
  spice_pullup pullup_7802(reg_iyh0_v, reg_iyh0_port_3);
  spice_pullup pullup_7803(reg_ixh0_v, reg_ixh0_port_3);
  spice_pullup pullup_7804(reg_d0_v, reg_d0_port_3);
  spice_pullup pullup_7805(reg_dd0_v, reg_dd0_port_3);
  spice_pullup pullup_7806(reg_h0_v, reg_h0_port_3);
  spice_pullup pullup_7807(reg_hh0_v, reg_hh0_port_3);
  spice_pullup pullup_7808(reg_b0_v, reg_b0_port_3);
  spice_pullup pullup_7809(reg_bb0_v, reg_bb0_port_3);
  spice_pullup pullup_7810(reg_aa0_v, reg_aa0_port_3);
  spice_pullup pullup_7811(reg_a0_v, reg_a0_port_3);
  spice_pullup pullup_7815(reg_pch1_v, reg_pch1_port_3);
  spice_pullup pullup_7816(reg_i1_v, reg_i1_port_3);
  spice_pullup pullup_7818(reg_w1_v, reg_w1_port_3);
  spice_pullup pullup_7819(reg_sph1_v, reg_sph1_port_3);
  spice_pullup pullup_7820(reg_iyh1_v, reg_iyh1_port_3);
  spice_pullup pullup_7821(reg_ixh1_v, reg_ixh1_port_3);
  spice_pullup pullup_7822(reg_d1_v, reg_d1_port_3);
  spice_pullup pullup_7823(reg_dd1_v, reg_dd1_port_3);
  spice_pullup pullup_7824(reg_h1_v, reg_h1_port_3);
  spice_pullup pullup_7825(reg_hh1_v, reg_hh1_port_3);
  spice_pullup pullup_7826(reg_b1_v, reg_b1_port_3);
  spice_pullup pullup_7827(reg_bb1_v, reg_bb1_port_3);
  spice_pullup pullup_7828(reg_aa1_v, reg_aa1_port_3);
  spice_pullup pullup_7829(reg_a1_v, reg_a1_port_3);
  spice_pullup pullup_7832(n_2306_v, n_2306_port_3);
  spice_pullup pullup_7833(n_2307_v, n_2307_port_3);
  spice_pullup pullup_7835(n_2308_v, n_2308_port_3);
  spice_pullup pullup_7836(n_2309_v, n_2309_port_3);
  spice_pullup pullup_7837(n_2310_v, n_2310_port_3);
  spice_pullup pullup_7838(n_2311_v, n_2311_port_3);
  spice_pullup pullup_7839(n_2312_v, n_2312_port_3);
  spice_pullup pullup_7840(n_2313_v, n_2313_port_3);
  spice_pullup pullup_7841(n_2314_v, n_2314_port_3);
  spice_pullup pullup_7842(n_2315_v, n_2315_port_3);
  spice_pullup pullup_7843(n_2316_v, n_2316_port_3);
  spice_pullup pullup_7844(n_2317_v, n_2317_port_3);
  spice_pullup pullup_7845(n_2318_v, n_2318_port_3);
  spice_pullup pullup_7846(n_2319_v, n_2319_port_3);
  spice_pullup pullup_7852(n_2344_v, n_2344_port_3);
  spice_pullup pullup_7853(n_2345_v, n_2345_port_3);
  spice_pullup pullup_7854(n_2346_v, n_2346_port_3);
  spice_pullup pullup_7855(n_2347_v, n_2347_port_3);
  spice_pullup pullup_7856(n_2348_v, n_2348_port_3);
  spice_pullup pullup_7857(n_2349_v, n_2349_port_3);
  spice_pullup pullup_7858(n_2350_v, n_2350_port_3);
  spice_pullup pullup_7859(n_2351_v, n_2351_port_3);
  spice_pullup pullup_7860(n_2352_v, n_2352_port_3);
  spice_pullup pullup_7861(n_2353_v, n_2353_port_3);
  spice_pullup pullup_7862(n_2354_v, n_2354_port_3);
  spice_pullup pullup_7863(n_2355_v, n_2355_port_3);
  spice_pullup pullup_7864(n_2356_v, n_2356_port_3);
  spice_pullup pullup_7865(n_2357_v, n_2357_port_3);
  spice_pullup pullup_7871(reg_pch2_v, reg_pch2_port_3);
  spice_pullup pullup_7872(reg_i2_v, reg_i2_port_3);
  spice_pullup pullup_7873(reg_w2_v, reg_w2_port_3);
  spice_pullup pullup_7874(reg_sph2_v, reg_sph2_port_3);
  spice_pullup pullup_7875(reg_iyh2_v, reg_iyh2_port_3);
  spice_pullup pullup_7876(reg_ixh2_v, reg_ixh2_port_3);
  spice_pullup pullup_7877(reg_d2_v, reg_d2_port_3);
  spice_pullup pullup_7878(reg_dd2_v, reg_dd2_port_3);
  spice_pullup pullup_7879(reg_h2_v, reg_h2_port_3);
  spice_pullup pullup_7880(reg_hh2_v, reg_hh2_port_3);
  spice_pullup pullup_7881(reg_b2_v, reg_b2_port_3);
  spice_pullup pullup_7882(reg_bb2_v, reg_bb2_port_3);
  spice_pullup pullup_7883(reg_aa2_v, reg_aa2_port_3);
  spice_pullup pullup_7884(reg_a2_v, reg_a2_port_3);
  spice_pullup pullup_7889(reg_pch3_v, reg_pch3_port_3);
  spice_pullup pullup_7890(reg_i3_v, reg_i3_port_3);
  spice_pullup pullup_7892(reg_w3_v, reg_w3_port_3);
  spice_pullup pullup_7893(reg_sph3_v, reg_sph3_port_3);
  spice_pullup pullup_7894(reg_iyh3_v, reg_iyh3_port_3);
  spice_pullup pullup_7895(reg_ixh3_v, reg_ixh3_port_3);
  spice_pullup pullup_7896(reg_d3_v, reg_d3_port_3);
  spice_pullup pullup_7897(reg_dd3_v, reg_dd3_port_3);
  spice_pullup pullup_7898(reg_h3_v, reg_h3_port_3);
  spice_pullup pullup_7899(reg_hh3_v, reg_hh3_port_3);
  spice_pullup pullup_7900(reg_b3_v, reg_b3_port_3);
  spice_pullup pullup_7901(reg_bb3_v, reg_bb3_port_3);
  spice_pullup pullup_7902(reg_aa3_v, reg_aa3_port_3);
  spice_pullup pullup_7903(reg_a3_v, reg_a3_port_3);
  spice_pullup pullup_7906(n_2429_v, n_2429_port_3);
  spice_pullup pullup_7907(n_2430_v, n_2430_port_3);
  spice_pullup pullup_7908(n_2431_v, n_2431_port_3);
  spice_pullup pullup_7909(n_2432_v, n_2432_port_3);
  spice_pullup pullup_7910(n_2433_v, n_2433_port_3);
  spice_pullup pullup_7911(n_2434_v, n_2434_port_3);
  spice_pullup pullup_7912(n_2435_v, n_2435_port_3);
  spice_pullup pullup_7913(n_2436_v, n_2436_port_3);
  spice_pullup pullup_7914(n_2437_v, n_2437_port_3);
  spice_pullup pullup_7915(n_2438_v, n_2438_port_3);
  spice_pullup pullup_7916(n_2439_v, n_2439_port_3);
  spice_pullup pullup_7917(n_2440_v, n_2440_port_3);
  spice_pullup pullup_7918(n_2441_v, n_2441_port_3);
  spice_pullup pullup_7919(n_2442_v, n_2442_port_3);
  spice_pullup pullup_7925(n_2450_v, n_2450_port_3);
  spice_pullup pullup_7926(n_2451_v, n_2451_port_3);
  spice_pullup pullup_7927(n_2452_v, n_2452_port_3);
  spice_pullup pullup_7928(n_2453_v, n_2453_port_3);
  spice_pullup pullup_7929(n_2454_v, n_2454_port_3);
  spice_pullup pullup_7930(n_2455_v, n_2455_port_3);
  spice_pullup pullup_7931(n_2456_v, n_2456_port_3);
  spice_pullup pullup_7932(n_2457_v, n_2457_port_3);
  spice_pullup pullup_7933(n_2458_v, n_2458_port_3);
  spice_pullup pullup_7934(n_2459_v, n_2459_port_3);
  spice_pullup pullup_7935(n_2460_v, n_2460_port_3);
  spice_pullup pullup_7936(n_2461_v, n_2461_port_3);
  spice_pullup pullup_7937(n_2462_v, n_2462_port_3);
  spice_pullup pullup_7938(n_2463_v, n_2463_port_3);
  spice_pullup pullup_7944(reg_pch4_v, reg_pch4_port_3);
  spice_pullup pullup_7945(reg_i4_v, reg_i4_port_3);
  spice_pullup pullup_7946(reg_w4_v, reg_w4_port_3);
  spice_pullup pullup_7947(reg_sph4_v, reg_sph4_port_3);
  spice_pullup pullup_7948(reg_iyh4_v, reg_iyh4_port_3);
  spice_pullup pullup_7949(reg_ixh4_v, reg_ixh4_port_3);
  spice_pullup pullup_7950(reg_d4_v, reg_d4_port_3);
  spice_pullup pullup_7951(reg_dd4_v, reg_dd4_port_3);
  spice_pullup pullup_7952(reg_h4_v, reg_h4_port_3);
  spice_pullup pullup_7953(reg_hh4_v, reg_hh4_port_3);
  spice_pullup pullup_7954(reg_b4_v, reg_b4_port_3);
  spice_pullup pullup_7955(reg_bb4_v, reg_bb4_port_3);
  spice_pullup pullup_7956(reg_aa4_v, reg_aa4_port_3);
  spice_pullup pullup_7957(reg_a4_v, reg_a4_port_3);
  spice_pullup pullup_7963(reg_pch5_v, reg_pch5_port_3);
  spice_pullup pullup_7964(reg_i5_v, reg_i5_port_3);
  spice_pullup pullup_7966(reg_w5_v, reg_w5_port_3);
  spice_pullup pullup_7967(reg_sph5_v, reg_sph5_port_3);
  spice_pullup pullup_7968(reg_iyh5_v, reg_iyh5_port_3);
  spice_pullup pullup_7969(reg_ixh5_v, reg_ixh5_port_3);
  spice_pullup pullup_7970(reg_d5_v, reg_d5_port_3);
  spice_pullup pullup_7971(reg_dd5_v, reg_dd5_port_3);
  spice_pullup pullup_7972(reg_h5_v, reg_h5_port_3);
  spice_pullup pullup_7973(reg_hh5_v, reg_hh5_port_3);
  spice_pullup pullup_7974(reg_b5_v, reg_b5_port_3);
  spice_pullup pullup_7975(reg_bb5_v, reg_bb5_port_3);
  spice_pullup pullup_7976(reg_aa5_v, reg_aa5_port_3);
  spice_pullup pullup_7977(reg_a5_v, reg_a5_port_3);
  spice_pullup pullup_7980(n_2539_v, n_2539_port_3);
  spice_pullup pullup_7981(n_2540_v, n_2540_port_3);
  spice_pullup pullup_7982(n_2541_v, n_2541_port_3);
  spice_pullup pullup_7983(n_2542_v, n_2542_port_3);
  spice_pullup pullup_7984(n_2543_v, n_2543_port_3);
  spice_pullup pullup_7985(n_2544_v, n_2544_port_3);
  spice_pullup pullup_7986(n_2545_v, n_2545_port_3);
  spice_pullup pullup_7987(n_2546_v, n_2546_port_3);
  spice_pullup pullup_7988(n_2547_v, n_2547_port_3);
  spice_pullup pullup_7989(n_2548_v, n_2548_port_3);
  spice_pullup pullup_7990(n_2549_v, n_2549_port_3);
  spice_pullup pullup_7991(n_2550_v, n_2550_port_3);
  spice_pullup pullup_7992(n_2551_v, n_2551_port_3);
  spice_pullup pullup_7993(n_2552_v, n_2552_port_3);
  spice_pullup pullup_8000(n_2573_v, n_2573_port_3);
  spice_pullup pullup_8001(n_2574_v, n_2574_port_3);
  spice_pullup pullup_8002(n_2575_v, n_2575_port_3);
  spice_pullup pullup_8003(n_2576_v, n_2576_port_3);
  spice_pullup pullup_8004(n_2577_v, n_2577_port_3);
  spice_pullup pullup_8005(n_2578_v, n_2578_port_3);
  spice_pullup pullup_8006(n_2579_v, n_2579_port_3);
  spice_pullup pullup_8007(n_2580_v, n_2580_port_3);
  spice_pullup pullup_8008(n_2581_v, n_2581_port_3);
  spice_pullup pullup_8009(n_2582_v, n_2582_port_3);
  spice_pullup pullup_8010(n_2583_v, n_2583_port_3);
  spice_pullup pullup_8011(n_2584_v, n_2584_port_3);
  spice_pullup pullup_8012(n_2585_v, n_2585_port_3);
  spice_pullup pullup_8013(n_2586_v, n_2586_port_3);
  spice_pullup pullup_8019(reg_pch6_v, reg_pch6_port_3);
  spice_pullup pullup_8020(reg_i6_v, reg_i6_port_3);
  spice_pullup pullup_8021(reg_w6_v, reg_w6_port_3);
  spice_pullup pullup_8022(reg_sph6_v, reg_sph6_port_3);
  spice_pullup pullup_8023(reg_iyh6_v, reg_iyh6_port_3);
  spice_pullup pullup_8024(reg_ixh6_v, reg_ixh6_port_3);
  spice_pullup pullup_8025(reg_d6_v, reg_d6_port_3);
  spice_pullup pullup_8026(reg_dd6_v, reg_dd6_port_3);
  spice_pullup pullup_8027(reg_h6_v, reg_h6_port_3);
  spice_pullup pullup_8028(reg_hh6_v, reg_hh6_port_3);
  spice_pullup pullup_8029(reg_b6_v, reg_b6_port_3);
  spice_pullup pullup_8030(reg_bb6_v, reg_bb6_port_3);
  spice_pullup pullup_8031(reg_aa6_v, reg_aa6_port_3);
  spice_pullup pullup_8032(reg_a6_v, reg_a6_port_3);
  spice_pullup pullup_8036(reg_pch7_v, reg_pch7_port_3);
  spice_pullup pullup_8037(reg_i7_v, reg_i7_port_3);
  spice_pullup pullup_8039(reg_w7_v, reg_w7_port_3);
  spice_pullup pullup_8040(reg_sph7_v, reg_sph7_port_3);
  spice_pullup pullup_8041(reg_iyh7_v, reg_iyh7_port_3);
  spice_pullup pullup_8042(reg_ixh7_v, reg_ixh7_port_3);
  spice_pullup pullup_8043(reg_d7_v, reg_d7_port_3);
  spice_pullup pullup_8044(reg_dd7_v, reg_dd7_port_3);
  spice_pullup pullup_8045(reg_h7_v, reg_h7_port_3);
  spice_pullup pullup_8046(reg_hh7_v, reg_hh7_port_3);
  spice_pullup pullup_8047(reg_b7_v, reg_b7_port_3);
  spice_pullup pullup_8048(reg_bb7_v, reg_bb7_port_3);
  spice_pullup pullup_8049(reg_aa7_v, reg_aa7_port_3);
  spice_pullup pullup_8050(reg_a7_v, reg_a7_port_3);
  spice_pullup pullup_8052(n_2643_v, n_2643_port_3);
  spice_pullup pullup_8053(n_2644_v, n_2644_port_3);
  spice_pullup pullup_8054(n_2645_v, n_2645_port_3);
  spice_pullup pullup_8055(n_2646_v, n_2646_port_3);
  spice_pullup pullup_8056(n_2647_v, n_2647_port_3);
  spice_pullup pullup_8057(n_2648_v, n_2648_port_3);
  spice_pullup pullup_8058(n_2649_v, n_2649_port_3);
  spice_pullup pullup_8059(n_2650_v, n_2650_port_3);
  spice_pullup pullup_8060(n_2651_v, n_2651_port_3);
  spice_pullup pullup_8061(n_2652_v, n_2652_port_3);
  spice_pullup pullup_8062(n_2653_v, n_2653_port_3);
  spice_pullup pullup_8063(n_2654_v, n_2654_port_3);
  spice_pullup pullup_8064(n_2655_v, n_2655_port_3);
  spice_pullup pullup_8065(n_2656_v, n_2656_port_3);
  spice_pullup pullup_8090(n_1043_v, n_1043_port_3);
  spice_pullup pullup_8098(n_1072_v, n_1072_port_5);
  spice_pullup pullup_8100(n_1095_v, n_1095_port_4);
  spice_pullup pullup_8101(n_1076_v, n_1076_port_5);
  spice_pullup pullup_8103(n_1077_v, n_1077_port_5);
  spice_pullup pullup_8109(n_1092_v, n_1092_port_3);
  spice_pullup pullup_8114(n_1079_v, n_1079_port_3);
  spice_pullup pullup_8131(n_1080_v, n_1080_port_4);
  spice_pullup pullup_8139(n_1126_v, n_1126_port_5);
  spice_pullup pullup_8140(n_1171_v, n_1171_port_4);
  spice_pullup pullup_8155(n_1204_v, n_1204_port_3);
  spice_pullup pullup_8169(n_1220_v, n_1220_port_6);
  spice_pullup pullup_8215(n_1327_v, n_1327_port_2);
  spice_pullup pullup_8259(n_1466_v, n_1466_port_3);
  spice_pullup pullup_8275(n_1498_v, n_1498_port_2);
  spice_pullup pullup_8318(n_1586_v, n_1586_port_4);
  spice_pullup pullup_8337(n_1590_v, n_1590_port_3);
  spice_pullup pullup_8389(n_1783_v, n_1783_port_4);

  spice_latch latch_10386(eclk,ereset, n_684_v, v(n_903_v), n_2322_v);
  spice_latch latch_10387(eclk,ereset, v(clk_v), n_1413_v, n_1414_v);
  spice_latch latch_10388(eclk,ereset, v(clk_v), m4_v, n_1192_v);
  spice_latch latch_10389(eclk,ereset, v(clk_v), n_1531_v, n_1547_v);
  spice_latch latch_10390(eclk,ereset, v(clk_v), n_1550_v, n_1560_v);
  spice_latch latch_10391(eclk,ereset, v(clk_v), n_1530_v, n_1562_v);
  spice_latch latch_10392(eclk,ereset, v(clk_v), n_1532_v, n_1563_v);
  spice_latch latch_10393(eclk,ereset, v(clk_v), n_1518_v, n_1555_v);
  spice_latch latch_10394(eclk,ereset, v(clk_v), n_1571_v, n_1559_v);
  spice_latch latch_10395(eclk,ereset, v(clk_v), n_1205_v, n_1200_v);
  spice_latch latch_10396(eclk,ereset, v(clk_v), n_1699_v, n_644_v);
  spice_latch latch_10397(eclk,ereset, v(clk_v), n_116_v, n_1101_v);
  spice_latch latch_10398(eclk,ereset, v(clk_v), n_1345_v, n_1343_v);
  spice_latch latch_10399(eclk,ereset, v(clk_v), n_1538_v, n_1567_v);
  spice_latch latch_10400(eclk,ereset, v(clk_v), n_1542_v, n_1568_v);
  spice_latch latch_10401(eclk,ereset, v(n_475_v), n_1491_v, n_471_v);
  spice_latch latch_10402(eclk,ereset, v(clk_v), n_1276_v, n_1244_v);
  spice_latch latch_10403(eclk,ereset, v(clk_v), n_152_v, n_1138_v);
  spice_latch latch_10404(eclk,ereset, v(clk_v), n_1588_v, n_1570_v);
  spice_latch latch_10405(eclk,ereset, v(clk_v), n_645_v, n_1780_v);
  spice_latch latch_10406(eclk,ereset, v(clk_v), n_1539_v, n_1569_v);
  spice_latch latch_10407(eclk,ereset, v(clk_v), n_1176_v, n_1158_v);
  spice_latch latch_10408(eclk,ereset, v(clk_v), m2_v, n_1258_v);
  spice_latch latch_10409(eclk,ereset, v(clk_v), n_495_v, n_1575_v);
  spice_latch latch_10410(eclk,ereset, v(clk_v), n_524_v, n_1549_v);
  spice_latch latch_10411(eclk,ereset, v(clk_v), n_1311_v, n_1329_v);
  spice_latch latch_10412(eclk,ereset, v(clk_v), n_298_v, n_1319_v);
  spice_latch latch_10413(eclk,ereset, v(clk_v), n_1322_v, n_1323_v);
  spice_latch latch_10414(eclk,ereset, v(clk_v), n_1304_v, n_1324_v);
  spice_latch latch_10415(eclk,ereset, v(clk_v), n_1479_v, n_1499_v);
  spice_latch latch_10416(eclk,ereset, v(clk_v), n_1544_v, n_1603_v);
  spice_latch latch_10417(eclk,ereset, v(clk_v), n_530_v, n_1604_v);
  spice_latch latch_10418(eclk,ereset, v(clk_v), n_1091_v, n_1102_v);
  spice_latch latch_10419(eclk,ereset, v(clk_v), n_1166_v, n_1122_v);
  spice_latch latch_10420(eclk,ereset, v(clk_v), n_1131_v, n_1114_v);
  spice_latch latch_10421(eclk,ereset, n_684_v, v(n_889_v), n_2443_v);
  spice_latch latch_10422(eclk,ereset, v(clk_v), n_1806_v, n_1724_v);
  spice_latch latch_10423(eclk,ereset, v(clk_v), n_1199_v, n_1160_v);
  spice_latch latch_10424(eclk,ereset, v(clk_v), n_1431_v, n_1433_v);
  spice_latch latch_10425(eclk,ereset, v(clk_v), n_426_v, n_1436_v);
  spice_latch latch_10426(eclk,ereset, v(clk_v), n_443_v, n_1435_v);
  spice_latch latch_10427(eclk,ereset, v(clk_v), n_438_v, n_1437_v);
  spice_latch latch_10428(eclk,ereset, v(clk_v), n_411_v, n_1438_v);
  spice_latch latch_10429(eclk,ereset, v(clk_v), n_63_v, n_1052_v);
  spice_latch latch_10430(eclk,ereset, v(clk_v), n_1283_v, n_1269_v);
  spice_latch latch_10431(eclk,ereset, v(clk_v), _t2_v, n_1222_v);
  spice_latch latch_10432(eclk,ereset, v(clk_v), n_1582_v, n_1597_v);
  spice_latch latch_10433(eclk,ereset, v(clk_v), m3_v, n_1124_v);
  spice_latch latch_10434(eclk,ereset, v(clk_v), n_99_v, n_1107_v);
  spice_latch latch_10435(eclk,ereset, v(clk_v), n_1206_v, n_1219_v);
  spice_latch latch_10436(eclk,ereset, v(clk_v), n_269_v, n_1321_v);
  spice_latch latch_10437(eclk,ereset, v(clk_v), n_549_v, n_1611_v);
  spice_latch latch_10438(eclk,ereset, v(clk_v), n_538_v, n_1613_v);
  spice_latch latch_10439(eclk,ereset, v(clk_v), n_95_v, n_1059_v);
  spice_latch latch_10440(eclk,ereset, n_684_v, n_943_v, n_2493_v);
  spice_latch latch_10441(eclk,ereset, v(clk_v), n_497_v, n_1602_v);
  spice_latch latch_10442(eclk,ereset, n_684_v, v(n_951_v), n_2474_v);
  spice_latch latch_10443(eclk,ereset, v(clk_v), n_558_v, n_1564_v);
  spice_latch latch_10444(eclk,ereset, v(clk_v), n_1294_v, n_1253_v);
  spice_latch latch_10445(eclk,ereset, v(clk_v), n_1208_v, n_1251_v);
  spice_latch latch_10446(eclk,ereset, v(clk_v), n_1281_v, n_1272_v);
  spice_latch latch_10447(eclk,ereset, v(clk_v), n_558_v, n_1610_v);
  spice_latch latch_10448(eclk,ereset, v(clk_v), n_1353_v, n_1356_v);
  spice_latch latch_10449(eclk,ereset, v(clk_v), n_1628_v, n_1614_v);
  spice_latch latch_10450(eclk,ereset, v(clk_v), n_454_v, n_1512_v);
  spice_latch latch_10451(eclk,ereset, v(clk_v), n_1224_v, n_1227_v);
  spice_latch latch_10452(eclk,ereset, v(clk_v), n_264_v, n_1331_v);
  spice_latch latch_10453(eclk,ereset, v(clk_v), n_548_v, n_559_v);
  spice_latch latch_10454(eclk,ereset, v(clk_v), n_66_v, n_1234_v);
  spice_latch latch_10455(eclk,ereset, v(clk_v), n_189_v, n_1240_v);
  spice_latch latch_10456(eclk,ereset, v(clk_v), n_531_v, n_1630_v);
  spice_latch latch_10457(eclk,ereset, v(clk_v), n_1694_v, n_1861_v);
  spice_latch latch_10458(eclk,ereset, v(clk_v), n_101_v, n_1342_v);
  spice_latch latch_10459(eclk,ereset, v(clk_v), n_758_v, n_1782_v);
  spice_latch latch_10460(eclk,ereset, v(clk_v), n_817_v, n_1810_v);
  spice_latch latch_10461(eclk,ereset, v(clk_v), _t3_v, n_1230_v);
  spice_latch latch_10462(eclk,ereset, n_684_v, v(n_937_v), n_2595_v);
  spice_latch latch_10463(eclk,ereset, n_684_v, n_844_v, n_2183_v);
  spice_latch latch_10464(eclk,ereset, v(clk_v), n_1573_v, n_1664_v);
  spice_latch latch_10465(eclk,ereset, n_684_v, v(n_852_v), n_2161_v);
  spice_latch latch_10466(eclk,ereset, v(clk_v), n_1648_v, n_1666_v);
  spice_latch latch_10467(eclk,ereset, v(clk_v), n_579_v, n_580_v);
  spice_latch latch_10468(eclk,ereset, n_684_v, v(n_545_v), n_1809_v);
  spice_latch latch_10469(eclk,ereset, v(clk_v), n_151_v, n_1159_v);
  spice_latch latch_10470(eclk,ereset, v(clk_v), n_1596_v, n_1652_v);
  spice_latch latch_10471(eclk,ereset, v(clk_v), n_564_v, n_1667_v);
  spice_latch latch_10472(eclk,ereset, v(clk_v), n_399_v, n_1398_v);
  spice_latch latch_10473(eclk,ereset, v(clk_v), n_1148_v, n_1134_v);
  spice_latch latch_10474(eclk,ereset, n_684_v, n_989_v, n_2657_v);
  spice_latch latch_10475(eclk,ereset, v(clk_v), n_527_v, n_1659_v);
  spice_latch latch_10476(eclk,ereset, n_684_v, v(n_995_v), n_2635_v);
  spice_latch latch_10477(eclk,ereset, v(clk_v), n_1662_v, n_1670_v);
  spice_latch latch_10478(eclk,ereset, v(clk_v), n_1546_v, n_1677_v);
  spice_latch latch_10479(eclk,ereset, v(clk_v), n_584_v, n_1663_v);
  spice_latch latch_10480(eclk,ereset, v(clk_v), n_1647_v, n_1675_v);
  spice_latch latch_10481(eclk,ereset, v(clk_v), n_1641_v, n_1676_v);
  spice_latch latch_10482(eclk,ereset, v(clk_v), n_1633_v, n_1681_v);
  spice_latch latch_10483(eclk,ereset, n_684_v, v(n_779_v), n_1864_v);
  spice_latch latch_10484(eclk,ereset, v(clk_v), n_1187_v, n_1174_v);
  spice_latch latch_10485(eclk,ereset, v(clk_v), n_1671_v, n_1669_v);
  spice_latch latch_10486(eclk,ereset, v(clk_v), n_1252_v, n_1261_v);
  spice_latch latch_10487(eclk,ereset, n_684_v, v(n_983_v), n_2694_v);
  spice_latch latch_10488(eclk,ereset, v(clk_v), n_1686_v, n_1660_v);
  spice_latch latch_10489(eclk,ereset, v(clk_v), n_1274_v, n_1235_v);
  spice_latch latch_10490(eclk,ereset, v(clk_v), n_593_v, n_1685_v);
  spice_latch latch_10491(eclk,ereset, v(clk_v), n_1085_v, n_1096_v);
  spice_latch latch_10492(eclk,ereset, v(clk_v), m1_v, n_1135_v);
  spice_latch latch_10493(eclk,ereset, v(clk_v), n_1690_v, n_1700_v);
  spice_latch latch_10494(eclk,ereset, v(clk_v), n_622_v, n_1704_v);
  spice_latch latch_10495(eclk,ereset, v(clk_v), n_1526_v, n_1527_v);
  spice_latch latch_10496(eclk,ereset, v(clk_v), n_187_v, n_1163_v);
  spice_latch latch_10497(eclk,ereset, v(clk_v), n_1291_v, n_1306_v);
  spice_latch latch_10498(eclk,ereset, v(clk_v), n_1275_v, n_1307_v);
  spice_latch latch_10499(eclk,ereset, v(clk_v), _t5_v, n_1157_v);
  spice_latch latch_10500(eclk,ereset, v(clk_v), n_1529_v, n_1535_v);
  spice_latch latch_10501(eclk,ereset, v(clk_v), n_1139_v, n_1162_v);
  spice_latch latch_10502(eclk,ereset, v(clk_v), n_540_v, n_1718_v);
  spice_latch latch_10503(eclk,ereset, n_684_v, v(n_837_v), n_2276_v);
  spice_latch latch_10504(eclk,ereset, v(clk_v), _t1_v, n_1183_v);
  spice_latch latch_10505(eclk,ereset, v(clk_v), n_1684_v, n_1720_v);
  spice_latch latch_10506(eclk,ereset, v(clk_v), n_1623_v, n_1721_v);
  spice_latch latch_10507(eclk,ereset, v(clk_v), n_500_v, n_1537_v);
  spice_latch latch_10508(eclk,ereset, v(clk_v), n_281_v, n_1416_v);
  spice_latch latch_10509(eclk,ereset, v(clk_v), n_1691_v, n_1726_v);
  spice_latch latch_10510(eclk,ereset, v(clk_v), n_1697_v, n_1729_v);
  spice_latch latch_10511(eclk,ereset, v(clk_v), n_1698_v, n_1734_v);
  spice_latch latch_10512(eclk,ereset, v(clk_v), n_1692_v, n_1735_v);
  spice_latch latch_10513(eclk,ereset, v(clk_v), _t4_v, n_1212_v);
  spice_latch latch_10514(eclk,ereset, v(clk_v), n_501_v, n_1543_v);
  spice_latch latch_10515(eclk,ereset, v(clk_v), n_621_v, n_1754_v);
  spice_latch latch_10516(eclk,ereset, n_684_v, n_896_v, n_2327_v);
  spice_latch latch_10517(eclk,ereset, (n_632_v&n_632_v), v(n_1701_v), n_1730_v);
  spice_latch latch_10518(eclk,ereset, (n_632_v&n_632_v), v(ex_dehl0_v), n_1731_v);
  spice_latch latch_10519(eclk,ereset, (v(clk_v)&n_608_v), v(n_769_v), n_1972_v);
  spice_latch latch_10520(eclk,ereset, (n_632_v&n_632_v), v(n_1702_v), n_1727_v);
  spice_latch latch_10521(eclk,ereset, (n_632_v&n_632_v), v(ex_dehl1_v), n_1728_v);
  spice_latch latch_10522(eclk,ereset, (n_624_v&n_624_v), v(ex_af_v), n_1767_v);
  spice_latch latch_10523(eclk,ereset, (n_624_v&n_624_v), v(n_633_v), n_1768_v);
  spice_latch latch_10524(eclk,ereset, (n_632_v&n_632_v), v(ex_bcdehl_v), n_1771_v);
  spice_latch latch_10525(eclk,ereset, (n_632_v&n_632_v), v(n_1773_v), n_1772_v);
  spice_latch latch_10526(eclk,ereset, (v(clk_v)&n_608_v), v(n_913_v), n_2394_v);
  spice_latch latch_10527(eclk,ereset, (v(clk_v)&n_608_v), v(n_929_v), n_2402_v);
  spice_latch latch_10528(eclk,ereset, (v(clk_v)&n_608_v), v(n_784_v), n_2065_v);
  spice_latch latch_10529(eclk,ereset, (n_436_v&v(clk_v)), n_691_v, n_1781_v);
  spice_latch latch_10530(eclk,ereset, (v(clk_v)&n_608_v), v(n_804_v), n_2068_v);
  spice_latch latch_10531(eclk,ereset, (v(clk_v)&n_608_v), v(n_948_v), n_2507_v);
  spice_latch latch_10532(eclk,ereset, (v(clk_v)&n_608_v), v(n_964_v), n_2513_v);
  spice_latch latch_10533(eclk,ereset, (v(clk_v)&n_608_v), v(n_707_v), n_1863_v);
  spice_latch latch_10534(eclk,ereset, (v(clk_v)&n_608_v), v(n_833_v), n_2159_v);
  spice_latch latch_10535(eclk,ereset, (v(clk_v)&n_747_v), v(n_728_v), n_1807_v);
  spice_latch latch_10536(eclk,ereset, (v(clk_v)&n_747_v), n_817_v, n_1831_v);
  spice_latch latch_10537(eclk,ereset, (v(clk_v)&n_608_v), v(n_857_v), n_2165_v);
  spice_latch latch_10538(eclk,ereset, (v(clk_v)&n_608_v), v(n_979_v), n_2614_v);
  spice_latch latch_10539(eclk,ereset, (v(clk_v)&n_608_v), v(n_722_v), n_1867_v);
  spice_latch latch_10540(eclk,ereset, (v(clk_v)&n_608_v), v(n_994_v), n_2619_v);
  spice_latch latch_10541(eclk,ereset, (v(clk_v)&n_608_v), v(n_879_v), n_2278_v);
  spice_latch latch_10542(eclk,ereset, (v(clk_v)&n_608_v), v(n_893_v), n_2282_v);
  spice_latch latch_10543(eclk,ereset, (v(clk_v)&n_608_v), v(n_744_v), n_1967_v);

  assign n_53_v = ~(v(_wait_v));
  assign n_63_v = ~((n_1049_v|v(n_1053_v)|n_74_v));
  assign n_74_v = ~((n_76_v|v(clk_v)|n_90_v));
  assign n_76_v = ~(n_1102_v);
  assign n_91_v = ~((n_1046_v|v(n_62_v)));
  assign n_102_v = ~(n_90_v);
  assign n_104_v = ~((v(n_75_v)|n_74_v|n_91_v));
  assign n_141_v = ~(n_186_v);
  assign n_151_v = ~((_t3_v|n_1173_v));
  assign n_153_v = ~((n_95_v|v(clk_v)|n_1200_v));
  assign n_154_v = ~(v(n_1184_v));
  assign n_158_v = ~(n_1151_v);
  assign n_167_v = ~(n_1177_v);
  assign n_174_v = ~(n_72_v);
  assign n_184_v = ~(((n_1233_v|n_194_v)|(n_233_v&m1_v)));
  assign n_186_v = ~(n_1244_v);
  assign n_193_v = ~(n_1253_v);
  assign n_198_v = ~((((n_95_v|m5_v)|(n_213_v&m4_v)|(m2_v&(n_203_v&n_1285_v)))|(m3_v&(n_287_v|(n_251_v&(n_1298_v|n_234_v))))));
  assign n_202_v = ~((n_295_v|n_309_v|n_311_v|n_340_v|n_301_v|n_345_v));
  assign n_203_v = ~(n_202_v);
  assign n_208_v = ~((m1_v&(n_1222_v&n_188_v)));
  assign n_211_v = ~((m1_v&(_t3_v|_t4_v)));
  assign n_212_v = ~(((n_232_v&n_1256_v)|(n_239_v&n_221_v)));
  assign n_213_v = ~(n_377_v);
  assign n_215_v = ~((n_256_v&n_235_v));
  assign n_217_v = ~(n_253_v);
  assign n_221_v = ~(n_232_v);
  assign n_224_v = ~(n_1324_v);
  assign n_233_v = ~((n_203_v|n_1337_v|n_232_v|n_1352_v));
  assign n_234_v = ~(n_402_v);
  assign n_235_v = ~(((_t4_v&(n_242_v&m1_v))|(_t5_v&n_243_v)));
  assign n_238_v = ~((n_264_v|n_269_v|n_298_v));
  assign n_239_v = ~((n_228_v|n_289_v|n_290_v|n_295_v|n_272_v|n_349_v|n_300_v|n_237_v|n_294_v|n_331_v|n_346_v));
  assign n_242_v = ~((n_270_v|n_228_v|n_336_v|n_288_v|n_315_v|n_334_v|n_325_v|n_324_v|n_340_v|n_300_v));
  assign n_243_v = ~((n_334_v|n_336_v));
  assign n_246_v = ~((n_1230_v&n_129_v));
  assign n_251_v = ~((n_318_v|n_325_v|n_324_v|n_302_v|n_363_v|n_339_v|n_342_v|n_292_v|n_343_v|n_344_v|n_347_v|n_303_v|n_270_v));
  assign n_252_v = ~(((n_217_v&m4_v)|(n_325_v&m3_v)|(n_324_v&m2_v)));
  assign n_253_v = ~((n_295_v|n_290_v));
  assign n_256_v = ~((_t6_v|(n_1351_v&_t3_v)|(n_372_v&_t4_v)));
  assign n_257_v = ~((n_262_v|n_220_v|n_330_v));
  assign n_260_v = ~(((m2_v|(n_1355_v&m5_v)|(n_257_v&m4_v))|(m3_v&(n_234_v|(n_329_v&n_194_v)))));
  assign n_261_v = ~((n_265_v|n_1347_v|n_1358_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_262_v = ~(n_432_v);
  assign n_287_v = ~((n_265_v|n_1364_v|n_1368_v|n_1377_v|n_247_v|n_1393_v));
  assign n_288_v = ~((n_267_v|n_374_v|n_1358_v|n_378_v|n_1371_v|n_1377_v|v(n_248_v)));
  assign n_289_v = ~((n_267_v|n_374_v|n_1358_v|n_1371_v|n_1377_v|v(n_248_v)));
  assign n_290_v = ~((n_265_v|n_1358_v|n_1364_v|n_1371_v|n_1373_v));
  assign n_291_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|v(n_248_v)|n_247_v|n_1390_v));
  assign n_292_v = ~((n_265_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1373_v));
  assign n_293_v = ~((n_265_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1373_v|v(n_248_v)));
  assign n_308_v = ~((n_192_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|n_385_v|n_247_v|n_1390_v));
  assign n_313_v = ~((n_267_v|n_374_v|n_375_v|n_378_v|n_1368_v|n_1373_v|n_1390_v));
  assign n_314_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|n_385_v|n_247_v|n_1393_v));
  assign n_315_v = ~((n_265_v|n_374_v|n_375_v|n_378_v|n_1371_v|n_1373_v|n_1390_v));
  assign n_316_v = ~((n_267_v|n_374_v|n_1358_v|n_1364_v|n_1371_v|n_1377_v|n_385_v|n_247_v|n_1393_v));
  assign n_317_v = ~((n_267_v|n_1347_v|n_375_v|n_1364_v|n_1368_v|n_1373_v|n_1390_v));
  assign n_318_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|v(n_248_v)|n_247_v|n_1393_v));
  assign n_319_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1368_v|n_1373_v|n_385_v));
  assign n_320_v = ~((n_265_v|n_1347_v|n_1358_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_324_v = ~((n_265_v|n_1347_v|n_375_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_325_v = ~((n_265_v|n_374_v|n_375_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_329_v = ~((n_251_v|n_220_v|n_234_v));
  assign n_332_v = ~((n_267_v|n_374_v|n_1358_v|n_1364_v|n_1371_v|n_1377_v|n_385_v|n_1386_v|n_1390_v));
  assign n_333_v = ~((n_267_v|n_374_v|n_1358_v|n_378_v|n_1371_v|n_1377_v|n_385_v|n_1386_v));
  assign n_334_v = ~((n_267_v|n_374_v|n_1358_v|n_1364_v|n_1371_v|n_1377_v|n_385_v|n_1386_v|n_1393_v));
  assign n_335_v = ~((n_267_v|n_374_v|n_1358_v|n_1364_v|n_1368_v|n_1373_v|v(n_248_v)));
  assign n_336_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1368_v|n_1373_v));
  assign n_337_v = ~((n_267_v|n_1347_v|n_375_v|n_1364_v|n_1368_v|n_1373_v|v(n_248_v)));
  assign n_338_v = ~((n_267_v|n_1347_v|n_375_v|n_378_v|n_1368_v|n_1373_v));
  assign n_339_v = ~((n_267_v|n_374_v|n_1358_v|n_378_v|n_1371_v|n_1377_v|n_385_v|n_247_v|n_1390_v));
  assign n_340_v = ~((n_267_v|n_1347_v|n_1358_v|n_1364_v|n_1368_v|n_1373_v|v(n_248_v)|n_1386_v|n_1390_v));
  assign n_341_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|v(n_248_v)|n_1386_v|n_1390_v));
  assign n_342_v = ~((n_267_v|n_1347_v|n_375_v|n_1364_v|n_1368_v|n_1373_v|n_247_v|n_1393_v));
  assign n_52_v = ~(v(_nmi_v));
  assign n_55_v = ~(n_1101_v);
  assign n_60_v = ~(n_52_v);
  assign n_79_v = ~((n_97_v|n_106_v|n_114_v));
  assign n_97_v = ~((n_106_v|n_114_v|n_1099_v));
  assign n_109_v = ~(((n_1083_v|n_112_v)|(n_1084_v&v(clk_v))));
  assign n_112_v = ~((n_1114_v|v(clk_v)|n_65_v));
  assign n_113_v = ~(((v(n_148_v)|v(n_150_v)|n_108_v)|(n_1116_v&n_122_v)));
  assign n_114_v = ~((n_106_v|n_1122_v|v(n_1095_v)));
  assign n_116_v = ~((v(n_148_v)|n_95_v));
  assign n_117_v = ~(n_123_v);
  assign n_121_v = ~(n_1138_v);
  assign n_125_v = ~((n_107_v|n_65_v));
  assign n_130_v = ~(((n_1100_v|n_108_v|n_135_v|n_95_v)|(n_1136_v&n_188_v)));
  assign n_135_v = ~(v(n_1171_v));
  assign n_145_v = ~((n_107_v|n_65_v|n_1185_v));
  assign n_152_v = ~((n_110_v|n_1115_v|n_160_v|n_95_v));
  assign n_156_v = ~(n_309_v);
  assign n_160_v = ~(n_238_v);
  assign n_164_v = ~(n_156_v);
  assign n_171_v = ~((n_1240_v|v(clk_v)));
  assign n_178_v = ~(n_1167_v);
  assign n_180_v = ~((v(clk_v)|n_1219_v));
  assign n_182_v = ~(((n_227_v&n_1188_v)|(n_142_v&(n_135_v|n_1237_v))));
  assign n_183_v = ~((v(clk_v)|n_135_v|n_1227_v));
  assign n_187_v = ~(((n_107_v|n_65_v)|(m1_v&(_t3_v|n_188_v))));
  assign n_189_v = ~((n_107_v&_t1_v));
  assign n_191_v = ~(v(n_181_v));
  assign n_200_v = ~(n_1264_v);
  assign n_201_v = ~((n_1255_v|n_1259_v));
  assign n_207_v = ~((n_1269_v|v(clk_v)));
  assign n_218_v = ~(n_1268_v);
  assign n_219_v = ~(n_1284_v);
  assign n_226_v = ~((n_1255_v|(n_1264_v&n_204_v)));
  assign n_227_v = ~((n_267_v|n_374_v|n_375_v|n_378_v|n_1371_v|n_1377_v));
  assign n_229_v = ~((n_1260_v|n_236_v));
  assign n_231_v = ~((n_245_v|n_191_v));
  assign n_236_v = ~(n_1215_v);
  assign n_237_v = ~((n_265_v|n_374_v|n_1358_v|n_378_v|n_1371_v|n_1373_v));
  assign n_245_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|n_1386_v|n_1393_v));
  assign n_249_v = ~((n_265_v|n_1347_v|n_375_v|n_378_v|n_1371_v|n_1373_v));
  assign n_255_v = ~((n_1329_v|v(clk_v)));
  assign n_258_v = ~((n_267_v|n_1347_v|n_375_v|n_378_v|n_1371_v|n_1373_v|v(n_248_v)|n_1386_v|n_1393_v));
  assign n_264_v = ~((n_267_v|n_374_v|n_1358_v|n_378_v|n_1371_v|n_1377_v|n_385_v|n_247_v|n_1393_v));
  assign n_266_v = ~((n_267_v|n_1347_v|n_375_v|n_378_v|n_1368_v|n_1377_v));
  assign n_268_v = ~((n_1325_v|n_385_v|n_1386_v|n_1393_v));
  assign n_269_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|n_385_v|n_247_v|n_1390_v));
  assign n_271_v = ~((n_265_v|n_374_v|n_375_v|n_378_v|n_1371_v|n_1373_v|n_247_v|n_1393_v));
  assign n_272_v = ~((n_265_v|n_1347_v|n_375_v|n_1364_v|n_1371_v|n_1373_v));
  assign n_273_v = ~((n_263_v|n_1368_v|n_1373_v));
  assign n_274_v = ~((n_263_v|n_1371_v|n_1373_v));
  assign n_275_v = ~((n_263_v|n_1371_v|n_1377_v));
  assign n_276_v = ~((n_267_v|n_374_v|n_1358_v|n_378_v|n_1368_v|n_1373_v));
  assign n_277_v = ~((n_1325_v|v(n_248_v)|n_1386_v|n_1390_v));
  assign n_278_v = ~((n_1325_v|n_385_v|n_1386_v|n_1390_v));
  assign n_279_v = ~((n_1325_v|n_385_v|n_247_v|n_1390_v));
  assign n_280_v = ~((n_267_v|n_374_v|n_375_v|n_378_v|n_1368_v|n_1373_v|n_385_v|n_247_v|n_1393_v));
  assign n_281_v = ~((n_1278_v|n_265_v|n_374_v|n_375_v|n_378_v|n_1371_v|n_1373_v|n_1386_v|n_1390_v));
  assign n_282_v = ~((n_1325_v|v(n_248_v)|n_247_v|n_1390_v));
  assign n_283_v = ~((n_1325_v|v(n_248_v)|n_247_v|n_1393_v));
  assign n_284_v = ~((n_1325_v|v(n_248_v)|n_1386_v|n_1393_v));
  assign n_285_v = ~((n_265_v|n_374_v|n_375_v|n_378_v|n_1371_v|n_1373_v|n_1386_v|n_1390_v));
  assign n_286_v = ~((n_1325_v|n_385_v|n_247_v|n_1393_v));
  assign n_294_v = ~((n_267_v|n_374_v|n_1358_v|n_1364_v|n_1371_v|n_1377_v|n_385_v|n_247_v|n_1390_v));
  assign n_295_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|n_1386_v|n_1390_v));
  assign n_296_v = ~((n_267_v|n_1347_v|n_1358_v|n_1364_v|n_1368_v|n_1373_v|n_385_v|n_247_v|n_1390_v));
  assign n_297_v = ~((n_192_v|n_267_v|n_1347_v|n_375_v|n_378_v|n_1368_v|n_1373_v|v(n_248_v)|n_1386_v|n_1393_v));
  assign n_298_v = ~((n_267_v|n_374_v|n_1358_v|n_378_v|n_1371_v|n_1377_v|n_385_v|n_1386_v));
  assign n_299_v = ~((n_267_v|n_1347_v|n_375_v|n_1364_v|n_1371_v|n_1377_v));
  assign n_300_v = ~((n_267_v|n_1347_v|n_1358_v|n_1364_v|n_1371_v|n_1377_v));
  assign n_301_v = ~((n_267_v|n_1347_v|n_1358_v|n_1364_v|n_1368_v|n_1373_v|n_385_v|n_1386_v|n_1390_v));
  assign n_302_v = ~((n_192_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|n_385_v|n_247_v|n_1390_v));
  assign n_303_v = ~((n_192_v|n_263_v));
  assign n_304_v = ~((n_258_v|n_267_v|n_1347_v|n_375_v|n_378_v|n_1371_v|n_1373_v));
  assign n_305_v = ~((n_258_v|n_267_v|n_1371_v|n_1373_v|v(n_248_v)|n_1386_v|n_1393_v));
  assign n_306_v = ~(n_263_v);
  assign n_307_v = ~((n_267_v|n_1358_v|n_378_v|n_1368_v|n_1373_v));
  assign n_309_v = ~((n_267_v|n_1347_v|n_375_v|n_378_v|n_1368_v|n_1373_v));
  assign n_310_v = ~((n_1305_v|n_219_v));
  assign n_311_v = ~((n_267_v|n_1347_v|n_375_v|n_378_v|n_1371_v|n_1377_v));
  assign n_312_v = ~((n_267_v|n_1368_v|n_1377_v));
  assign n_321_v = ~((n_267_v|n_374_v|n_375_v|n_378_v|n_1368_v|n_1373_v|n_385_v|n_1386_v|n_1393_v));
  assign n_322_v = ~((n_265_v|n_375_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_323_v = ~((n_265_v|n_374_v|n_1358_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_331_v = ~((n_267_v|n_1347_v|n_375_v|n_1364_v|n_1368_v|n_1373_v|n_1390_v));
  assign n_343_v = ~((n_267_v|n_1347_v|n_375_v|n_1364_v|n_1368_v|n_1373_v|n_1386_v|n_1393_v));
  assign n_344_v = ~((n_267_v|n_1347_v|n_1358_v|n_378_v|n_1371_v|n_1377_v));
  assign n_345_v = ~((n_267_v|n_1347_v|n_1358_v|n_1364_v|n_1368_v|n_1373_v|n_1393_v));
  assign n_346_v = ~((n_267_v|n_1347_v|n_375_v|n_378_v|n_1368_v|n_1373_v|v(n_248_v)|n_1386_v|n_1393_v));
  assign n_347_v = ~((n_267_v|n_1358_v|n_378_v|n_1368_v|n_1373_v|v(n_248_v)|n_1386_v|n_1393_v));
  assign n_348_v = ~((n_267_v|n_1371_v|n_1373_v));
  assign n_349_v = ~((n_267_v|n_374_v|n_1358_v|n_1364_v|n_1368_v|n_1373_v|n_385_v));
  assign n_350_v = ~((n_267_v|n_374_v|n_375_v|n_378_v|n_1368_v|n_1373_v|n_1390_v));
  assign n_351_v = ~((n_263_v|n_1368_v|n_1377_v));
  assign n_352_v = ~((n_267_v|n_374_v|n_375_v|n_378_v|n_1368_v|n_1373_v|v(n_248_v)|n_247_v|n_1393_v));
  assign n_353_v = ~((n_267_v|n_1347_v|n_1358_v|n_1364_v|n_1368_v|n_1373_v|v(n_248_v)|n_1386_v|n_1390_v));
  assign n_354_v = ~((n_267_v|n_374_v|n_375_v|n_378_v|n_1368_v|n_1373_v|v(n_248_v)|n_1386_v|n_1393_v));
  assign n_355_v = ~((n_267_v|n_374_v|n_375_v|n_1364_v|n_1371_v|n_1377_v|n_1386_v|n_1390_v));
  assign n_356_v = ~((n_263_v|n_1347_v|n_375_v|n_378_v));
  assign n_357_v = ~(n_1348_v);
  assign n_360_v = ~((n_325_v|n_324_v|n_340_v|n_299_v|n_301_v|n_345_v|n_320_v|n_364_v|n_339_v|n_335_v|n_318_v|n_363_v|n_291_v|n_342_v|n_292_v|n_343_v|n_344_v|n_270_v));
  assign n_361_v = ~((n_265_v|n_374_v|n_1358_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_363_v = ~((n_265_v|n_374_v|n_375_v|n_378_v|n_1371_v|n_1373_v|n_247_v|n_1393_v));
  assign n_364_v = ~((n_265_v|n_374_v|n_1358_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_365_v = ~((n_265_v|n_374_v|n_375_v|n_378_v|n_1371_v|n_1373_v|n_1390_v));
  assign n_372_v = ~((n_1361_v|n_262_v));
  assign n_377_v = ~((n_363_v|n_320_v|n_364_v|n_325_v|n_324_v|n_290_v|n_331_v|n_295_v|n_343_v|n_346_v|n_305_v|n_266_v|n_304_v|n_274_v));
  assign n_381_v = ~((v(n_384_v)|(v(n_359_v)&n_78_v)));
  assign n_386_v = ~((n_389_v|n_65_v));
  assign n_389_v = ~(((n_270_v&m2_v)|(n_387_v&m4_v)|(m5_v&(n_387_v|n_220_v))|(m3_v&(n_262_v|n_270_v))));
  assign n_390_v = ~((_t1_v|(m1_v&_t3_v)));
  assign n_391_v = ~(n_1444_v);
  assign n_394_v = ~((n_1389_v|n_318_v));
  assign n_396_v = ~(((n_1396_v&(m5_v|m4_v))|(n_1399_v&m3_v)));
  assign n_398_v = ~((n_316_v|n_228_v|n_339_v|n_340_v|n_291_v|n_294_v|n_344_v|n_299_v|n_300_v|n_237_v|n_301_v|n_345_v|n_270_v));
  assign n_399_v = ~(((n_334_v&_t4_v)|(_t3_v&(n_318_v&m5_v))));
  assign n_401_v = ~(n_422_v);
  assign n_402_v = ~((n_335_v|n_291_v|n_342_v|n_292_v|n_343_v|n_299_v|n_270_v|n_325_v|n_324_v));
  assign n_407_v = ~(((_t4_v&(n_410_v&m1_v))|(_t3_v&(n_394_v&m3_v))|((_t1_v|_t3_v)&(n_262_v&m4_v))));
  assign n_410_v = ~((n_429_v&n_1412_v));
  assign n_416_v = ~((n_434_v|n_361_v|n_363_v));
  assign n_417_v = ~((n_348_v|n_306_v|n_311_v|n_312_v|n_307_v));
  assign n_419_v = ~(n_262_v);
  assign n_420_v = ~((n_336_v|n_334_v|n_318_v|n_337_v|n_288_v|n_339_v|n_363_v|n_341_v|n_344_v|n_293_v|n_362_v|n_346_v|n_305_v|n_228_v));
  assign n_422_v = ~((n_339_v|n_291_v|n_342_v|n_292_v|n_335_v|n_297_v|n_343_v|n_344_v|n_299_v|n_302_v|n_303_v));
  assign n_424_v = ~((n_318_v|n_289_v|n_339_v|n_294_v|n_300_v|n_237_v|n_228_v|n_344_v));
  assign n_429_v = ~((n_319_v|n_288_v));
  assign n_430_v = ~((n_340_v|n_301_v|n_345_v));
  assign n_432_v = ~((n_320_v|n_364_v|n_325_v|n_324_v));
  assign n_433_v = ~((n_339_v|n_344_v));
  assign n_434_v = ~((n_262_v|n_1502_v));
  assign n_435_v = ~((n_340_v|n_290_v|n_324_v|n_325_v));
  assign n_440_v = ~((((m1_v&_t3_v)|((n_270_v|n_387_v)&(_t5_v&m1_v)))|(_t2_v&((n_262_v&m3_v)|(m5_v&(n_395_v&n_456_v))))));
  assign n_441_v = ~((n_334_v|n_316_v|n_363_v|n_320_v|n_364_v|n_232_v));
  assign n_442_v = ~((n_313_v|n_340_v|n_325_v|n_324_v));
  assign n_446_v = ~((v(n_248_v)|n_467_v));
  assign n_453_v = ~(((m1_v|m3_v)|(n_1425_v&m2_v)));
  assign n_454_v = ~(((n_1432_v|n_465_v|n_1481_v)|(n_1476_v&(n_101_v|n_1449_v))));
  assign n_455_v = ~(n_433_v);
  assign n_457_v = ~(((n_478_v|n_1458_v|n_335_v|n_289_v|n_395_v)|(v(n_248_v)&n_1421_v)));
  assign n_459_v = ~(n_430_v);
  assign n_461_v = ~(((m1_v&_t4_v)|(_t2_v&(m1_v|(n_395_v&m3_v)))|(_t3_v&(m5_v|(n_262_v&m3_v)))));
  assign n_464_v = ~(n_442_v);
  assign n_466_v = ~((n_192_v|n_1448_v));
  assign n_467_v = ~((n_342_v|n_292_v));
  assign n_468_v = ~(n_427_v);
  assign n_470_v = ~((n_268_v|n_400_v));
  assign n_472_v = ~(((_t4_v&(n_262_v&m4_v))|((n_455_v|n_228_v)&(_t1_v&(m5_v|m4_v)))));
  assign n_473_v = ~((n_391_v&m3_v));
  assign n_477_v = ~(((_t1_v&(n_270_v&(m3_v|m2_v)))|(n_459_v&((_t2_v&m2_v)|(m3_v&_t3_v)))));
  assign n_478_v = ~(n_445_v);
  assign n_482_v = ~((n_477_v&n_472_v));
  assign n_483_v = ~((n_1477_v&n_422_v));
  assign n_489_v = ~((n_110_v|(n_490_v&(n_1508_v|n_1509_v))));
  assign n_490_v = ~(((n_401_v&m2_v)|(n_483_v&m1_v)|(n_262_v&m3_v)));
  assign n_492_v = ~((n_478_v|n_1470_v));
  assign n_493_v = ~((n_95_v|(_t1_v&(m1_v|(n_483_v&m2_v)|(n_401_v&m3_v)))));
  assign n_495_v = ~((n_465_v|n_489_v|n_482_v));
  assign n_497_v = ~((n_465_v|n_489_v));
  assign n_362_v = ~((n_265_v|n_374_v|n_1358_v|n_1364_v|n_1371_v|n_1373_v));
  assign n_366_v = ~((n_265_v|n_374_v|n_375_v|n_378_v|n_1371_v|n_1373_v|n_247_v|n_1390_v));
  assign n_367_v = ~((n_265_v|n_1347_v|n_1358_v|n_1364_v|n_1371_v|n_1373_v));
  assign n_368_v = ~((n_265_v|n_1347_v|n_1358_v|n_378_v|n_1371_v|n_1373_v));
  assign n_369_v = ~((n_265_v|n_1347_v|n_1358_v|n_1364_v|n_1368_v|n_1377_v|n_1393_v));
  assign n_373_v = ~(n_1359_v);
  assign n_376_v = ~(n_1365_v);
  assign n_379_v = ~(n_1369_v);
  assign n_382_v = ~(n_1374_v);
  assign n_388_v = ~(n_1379_v);
  assign n_392_v = ~(n_1387_v);
  assign n_397_v = ~(n_1394_v);
  assign n_400_v = ~((n_271_v|n_280_v|n_368_v|n_285_v|n_311_v|n_312_v|n_350_v|n_352_v));
  assign n_403_v = ~((n_348_v|n_367_v|n_309_v|n_311_v|n_312_v|n_273_v|n_350_v|n_352_v|n_285_v));
  assign n_404_v = ~((n_311_v|n_312_v|n_307_v|n_367_v|n_272_v|n_349_v|n_273_v|n_274_v|n_321_v|n_322_v|n_354_v|n_323_v|n_369_v));
  assign n_405_v = ~((n_228_v|n_348_v|n_309_v|n_280_v|n_368_v|n_285_v|n_367_v|n_273_v|n_350_v));
  assign n_409_v = ~((n_368_v|n_272_v|n_349_v|n_268_v|n_277_v|n_278_v|n_279_v|n_282_v|n_284_v|n_286_v));
  assign n_411_v = ~((n_307_v|n_272_v|n_268_v|n_277_v|n_278_v|n_279_v|n_368_v|n_282_v|n_285_v));
  assign n_413_v = ~((n_280_v|n_368_v|n_351_v|n_276_v|n_268_v|n_277_v|n_278_v|n_353_v|n_322_v|n_323_v));
  assign n_415_v = ~((n_285_v|n_271_v|n_311_v|n_312_v|n_307_v|n_273_v|n_274_v|n_352_v|n_368_v|n_353_v|n_322_v|n_323_v|n_367_v|n_272_v));
  assign n_421_v = ~((n_307_v|n_280_v|n_283_v|n_274_v|n_353_v|n_322_v));
  assign n_423_v = ~((n_272_v|n_278_v|n_279_v|n_321_v));
  assign n_425_v = ~((n_266_v|n_347_v|n_303_v|n_356_v|n_304_v|n_302_v|n_346_v|n_305_v));
  assign n_426_v = ~((n_275_v|n_284_v|n_286_v));
  assign n_427_v = ~((n_351_v|n_275_v|n_348_v|n_309_v|n_307_v|n_367_v|n_273_v));
  assign n_428_v = ~((n_283_v|n_321_v|n_354_v));
  assign n_431_v = ~((n_301_v|n_345_v|n_306_v|n_307_v|n_353_v|n_322_v));
  assign n_437_v = ~((n_306_v|n_312_v));
  assign n_438_v = ~((n_275_v|n_284_v));
  assign n_439_v = ~((n_321_v|n_322_v|n_354_v|n_323_v|n_369_v));
  assign n_443_v = ~((n_283_v|n_274_v|n_351_v));
  assign n_444_v = ~((n_353_v|n_322_v));
  assign n_445_v = ~((n_331_v|n_295_v|n_343_v));
  assign n_447_v = ~(n_450_v);
  assign n_448_v = ~((n_353_v|n_322_v|n_323_v));
  assign n_449_v = ~(v(n_248_v));
  assign n_450_v = ~((n_437_v&(n_1424_v|_t2_v)));
  assign n_458_v = ~((n_322_v|n_439_v));
  assign n_460_v = ~((n_413_v&n_1443_v));
  assign n_462_v = ~((n_345_v|n_1393_v));
  assign n_463_v = ~(n_1454_v);
  assign n_469_v = ~((n_425_v|n_192_v));
  assign n_487_v = ~(n_82_v);
  assign n_488_v = ~(n_457_v);
  assign n_491_v = ~(n_1453_v);
  assign n_496_v = ~(((_t3_v&(n_228_v&m5_v))|(_t2_v&(n_270_v&m3_v))|(_t1_v&(n_355_v&m2_v))));
  assign n_498_v = ~(((n_558_v|(_t5_v&(n_270_v&m1_v))|(_t2_v&(m2_v&(n_220_v|n_469_v)))|(_t3_v&(n_220_v&(m3_v|m4_v))))|(_t4_v&((n_330_v&m4_v)|(m1_v&(n_220_v|n_330_v))))));
  assign n_504_v = ~(n_482_v);
  assign n_505_v = ~((((_t1_v&(n_478_v&m4_v))|(_t4_v&(n_313_v&m1_v))|(_t2_v&(n_470_v&m1_v)))|((n_478_v&n_456_v)&(m4_v&_t3_v))));
  assign n_506_v = ~((((_t3_v&(n_330_v&(m4_v|m5_v)))|(_t2_v&(n_1503_v&m2_v)))|(_t4_v&((n_330_v&m4_v)|(n_363_v&m3_v)))));
  assign n_507_v = ~(((_t2_v&(n_324_v&m3_v))|(_t5_v&(n_325_v&m1_v))|((n_324_v|n_338_v)&(_t3_v&m2_v))|((n_330_v|n_1490_v)&(_t4_v&m1_v))));
  assign n_508_v = ~((((_t1_v&(n_1489_v&m2_v))|(_t5_v&(n_324_v&m1_v)))|(_t3_v&((n_262_v&m3_v)|(n_325_v&m2_v)))|(_t4_v&((n_262_v&m3_v)|(n_1489_v&m1_v)))));
  assign n_510_v = ~(((_t3_v&(n_335_v&(m3_v|m2_v)))|((_t5_v|_t4_v)&(m5_v|(m1_v&(n_317_v|n_336_v))))));
  assign n_511_v = ~((n_466_v&((_t2_v&m2_v)|(m3_v&_t3_v))));
  assign n_512_v = ~(((_t3_v&(n_478_v&m4_v))|(_t5_v&(n_220_v&m3_v))|(_t2_v&(n_470_v&m1_v))));
  assign n_513_v = ~(((_t2_v&(n_270_v&m2_v))|((_t5_v|_t4_v)&((n_395_v|n_270_v)&(m3_v|m1_v)))));
  assign n_514_v = ~(n_1781_v);
  assign n_518_v = ~((_t2_v&(n_468_v&m1_v)));
  assign n_519_v = ~((n_332_v&n_535_v));
  assign n_520_v = ~((n_517_v|(n_502_v&n_1522_v)|(v(n_1590_v)&n_1548_v)));
  assign n_521_v = ~((v(clk_v)|n_1551_v));
  assign n_522_v = ~(n_511_v);
  assign n_529_v = ~((n_522_v|n_536_v|n_1578_v|n_558_v|n_1580_v|n_1584_v|n_1605_v));
  assign n_531_v = ~((n_511_v&(n_1583_v|n_581_v)));
  assign n_532_v = ~(n_1561_v);
  assign n_534_v = ~((n_314_v&n_535_v));
  assign n_535_v = ~(n_1560_v);
  assign n_536_v = ~((n_513_v&n_1552_v));
  assign n_537_v = ~((_t4_v&(n_365_v&m1_v)));
  assign n_547_v = ~((m1_v&_t3_v));
  assign n_555_v = ~((n_1576_v|n_592_v|n_1616_v));
  assign n_556_v = ~((n_567_v&(n_537_v|n_484_v)));
  assign n_563_v = ~(n_484_v);
  assign n_564_v = ~((n_508_v&(n_555_v|n_565_v)));
  assign n_565_v = ~((n_548_v&n_484_v));
  assign n_566_v = ~((n_479_v|(n_567_v&n_518_v)));
  assign n_567_v = ~(((_t4_v&(n_1465_v&m1_v))|((n_290_v|n_1463_v)&(_t1_v&m4_v))));
  assign n_568_v = ~((n_548_v|n_484_v));
  assign n_572_v = ~((n_548_v|n_484_v));
  assign n_571_v = ~(n_549_v);
  assign n_577_v = ~(n_1614_v);
  assign n_578_v = ~(n_1666_v);
  assign n_579_v = ~((n_536_v|(n_1643_v&n_592_v)));
  assign n_581_v = ~((n_1578_v|(n_1646_v&(n_1636_v|n_592_v))));
  assign n_584_v = ~(((n_1605_v|n_558_v)|(n_572_v&(n_1576_v|n_566_v))));
  assign n_585_v = ~((n_518_v&(n_537_v|n_1608_v)));
  assign n_591_v = ~(n_1640_v);
  assign n_592_v = ~((n_1541_v&n_510_v));
  assign n_593_v = ~((n_581_v|n_1474_v));
  assign n_601_v = ~(n_1664_v);
  assign n_606_v = ~(n_1703_v);
  assign ex_dehl_combined_v = ~(((v(ex_dehl1_v)&n_634_v)|(v(ex_dehl0_v)&n_640_v)));
  assign n_628_v = ~((n_519_v&n_534_v));
  assign n_630_v = ~(n_600_v);
  assign n_632_v = ~((n_628_v|v(clk_v)));
  assign n_640_v = ~(n_634_v);
  assign n_655_v = ~((v(clk_v)|n_599_v));
  assign n_656_v = ~((v(clk_v)|n_602_v));
  assign n_659_v = ~((v(clk_v)|n_1738_v));
  assign n_660_v = ~((v(clk_v)|n_1739_v));
  assign n_663_v = ~((v(clk_v)|n_1740_v));
  assign n_664_v = ~((v(clk_v)|n_1741_v));
  assign n_667_v = ~((v(clk_v)|n_1742_v));
  assign n_668_v = ~((v(clk_v)|n_1743_v));
  assign n_671_v = ~((v(clk_v)|n_1744_v));
  assign n_672_v = ~((v(clk_v)|n_1745_v));
  assign n_675_v = ~((v(clk_v)|n_1746_v));
  assign n_676_v = ~((v(clk_v)|n_1747_v));
  assign n_685_v = ~(n_577_v);
  assign n_690_v = ~((v(n_617_v)|n_406_v|v(n_709_v)|v(n_721_v)|v(n_746_v)|v(n_763_v)|v(n_787_v)|v(n_802_v)|v(n_835_v)));
  assign n_691_v = ~((n_1777_v|n_1886_v|n_1914_v|n_1992_v|n_2018_v|n_2088_v|n_2118_v|n_2187_v|n_2225_v|n_2301_v|n_2343_v|n_2422_v|n_2449_v|n_2534_v|n_2572_v|n_2660_v));
  assign n_694_v = ~(n_406_v);
  assign n_705_v = ~(n_706_v);
  assign n_706_v = ~((n_607_v|n_1863_v));
  assign n_710_v = ~((n_406_v|v(n_709_v)|v(n_721_v)));
  assign n_718_v = ~(n_725_v);
  assign n_725_v = ~((n_1867_v|n_607_v));
  assign n_730_v = ~(n_710_v);
  assign n_742_v = ~(n_743_v);
  assign n_743_v = ~((n_607_v|n_1967_v));
  assign n_748_v = ~((n_730_v|v(n_746_v)|v(n_763_v)));
  assign n_760_v = ~(n_771_v);
  assign n_771_v = ~((n_1972_v|n_607_v));
  assign n_773_v = ~(n_748_v);
  assign n_778_v = ~(v(n_2116_v));
  assign n_781_v = ~(n_782_v);
  assign n_782_v = ~((n_607_v|n_2065_v));
  assign n_789_v = ~((n_773_v|v(n_787_v)|v(n_802_v)));
  assign n_800_v = ~(n_805_v);
  assign n_805_v = ~((n_2068_v|n_607_v));
  assign n_811_v = ~(n_690_v);
  assign n_814_v = ~(n_815_v);
  assign n_815_v = ~((n_607_v|n_2159_v));
  assign n_842_v = ~((n_811_v|v(n_856_v)|v(n_881_v)|v(n_892_v)|v(n_915_v)|v(n_928_v)));
  assign n_851_v = ~(n_858_v);
  assign n_854_v = ~((n_811_v|v(n_856_v)|v(n_881_v)));
  assign n_858_v = ~((n_2165_v|n_607_v));
  assign n_499_v = ~(((m3_v&_t5_v)|(_t1_v&(n_220_v&(m2_v|m5_v)))|(_t3_v&(n_330_v&m5_v))|((n_470_v|n_468_v)&(m1_v&_t2_v))));
  assign n_500_v = ~((((_t1_v&(n_1483_v&m2_v))|(_t3_v&(n_330_v&m4_v)))|(_t2_v&((n_323_v&m3_v)|(n_448_v&m1_v)))));
  assign n_501_v = ~(n_1519_v);
  assign n_503_v = ~(((n_345_v&m2_v)|(n_1488_v&m3_v)|(n_300_v&m1_v)));
  assign n_515_v = ~(n_737_v);
  assign n_516_v = ~((((_t3_v|_t1_v)&(n_270_v&m2_v))|(_t4_v&(m4_v|(n_464_v&m1_v)))));
  assign n_517_v = ~((n_1566_v|n_1528_v));
  assign n_523_v = ~(((_t1_v&(n_488_v&m5_v))|(_t4_v&(n_491_v&m1_v))));
  assign n_524_v = ~(n_1517_v);
  assign n_527_v = ~((n_1571_v|n_540_v|n_1540_v|n_1542_v));
  assign n_530_v = ~(((n_1539_v|n_1545_v)|(n_524_v&n_463_v)));
  assign n_533_v = ~(((m2_v&_t2_v)|(_t1_v&((n_491_v&m4_v)|(n_270_v&m3_v)))));
  assign n_538_v = ~(((n_558_v|n_539_v)|(n_556_v&(n_479_v|n_568_v))));
  assign n_539_v = ~((n_1558_v&n_516_v));
  assign n_540_v = ~((n_499_v&n_1689_v));
  assign n_542_v = ~(n_1537_v);
  assign n_543_v = ~((n_1564_v&n_1565_v));
  assign n_550_v = ~(n_1611_v);
  assign n_554_v = ~((n_568_v|n_479_v));
  assign n_561_v = ~((n_524_v|n_501_v|n_1596_v));
  assign n_569_v = ~(n_479_v);
  assign n_573_v = ~(n_1613_v);
  assign n_582_v = ~((n_1494_v&n_612_v));
  assign n_583_v = ~(n_1604_v);
  assign n_594_v = ~(n_1446_v);
  assign n_598_v = ~(n_1669_v);
  assign n_605_v = ~(n_462_v);
  assign n_609_v = ~(n_605_v);
  assign n_610_v = ~(n_1670_v);
  assign n_611_v = ~((v(clk_v)|n_750_v));
  assign n_619_v = ~(n_1677_v);
  assign n_620_v = ~(n_1687_v);
  assign n_621_v = ~((_t2_v&(n_310_v&m4_v)));
  assign n_622_v = ~(((n_1459_v&n_612_v)|(_t4_v&(n_330_v&m4_v))|(_t3_v&(n_220_v&m3_v))));
  assign n_623_v = ~((n_1486_v&n_612_v));
  assign n_624_v = ~((n_619_v|v(clk_v)));
  assign n_635_v = ~(n_1732_v);
  assign n_636_v = ~((n_1688_v|v(clk_v)|n_638_v));
  assign n_637_v = ~((n_623_v|v(clk_v)));
  assign n_638_v = ~((n_1683_v&(n_1672_v|n_1536_v)));
  assign n_639_v = ~((n_1765_v|v(clk_v)));
  assign n_642_v = ~((n_1750_v|(n_635_v&n_1752_v)));
  assign n_645_v = ~((_t2_v&(n_1447_v&m1_v)));
  assign n_648_v = ~((n_638_v|v(clk_v)));
  assign n_649_v = ~(n_1720_v);
  assign n_650_v = ~((v(clk_v)|n_724_v));
  assign n_653_v = ~((v(clk_v)|n_620_v));
  assign n_679_v = ~((v(clk_v)|n_606_v));
  assign n_682_v = ~((n_1778_v&n_1760_v));
  assign n_683_v = ~(n_1423_v);
  assign n_686_v = ~(v(n_647_v));
  assign n_688_v = ~(((v(n_716_v)&n_1749_v)|(v(n_526_v)&n_1750_v)|(v(n_525_v)&n_1751_v)|(v(n_545_v)&n_1752_v)));
  assign n_698_v = ~(n_1807_v);
  assign n_699_v = ~(n_827_v);
  assign n_704_v = ~(v(n_545_v));
  assign n_711_v = ~(v(n_697_v));
  assign n_712_v = ~((n_1693_v|v(clk_v)));
  assign n_717_v = ~((n_1859_v&n_795_v));
  assign n_719_v = ~(v(n_528_v));
  assign n_720_v = ~(n_618_v);
  assign n_724_v = ~((n_1857_v&n_618_v));
  assign n_727_v = ~(v(n_728_v));
  assign n_736_v = ~((n_717_v|v(clk_v)));
  assign n_737_v = ~(n_1839_v);
  assign n_741_v = ~(v(n_526_v));
  assign n_756_v = ~((n_1723_v|(n_612_v&(n_220_v&n_1622_v))));
  assign n_758_v = ~(n_764_v);
  assign n_759_v = ~(n_818_v);
  assign n_761_v = ~(v(n_770_v));
  assign n_762_v = ~((n_2662_v&(n_2332_v|n_2498_v)));
  assign n_764_v = ~(v(n_726_v));
  assign n_765_v = ~(n_1858_v);
  assign n_766_v = ~(n_711_v);
  assign n_768_v = ~(n_729_v);
  assign n_780_v = ~(v(n_779_v));
  assign n_786_v = ~(n_751_v);
  assign n_788_v = ~(n_786_v);
  assign n_801_v = ~(v(n_790_v));
  assign n_812_v = ~(v(n_716_v));
  assign n_818_v = ~((n_2061_v|n_2184_v|v(n_2211_v)|n_2328_v|v(n_2338_v)|n_2494_v|v(n_2504_v)|n_2658_v|v(n_816_v)));
  assign n_819_v = ~((n_2682_v&((n_2390_v|n_2556_v)|(n_862_v&n_2226_v))));
  assign n_825_v = ~((n_1436_v|m6_v));
  assign n_826_v = ~((n_1435_v|m6_v));
  assign n_828_v = ~((n_1437_v|m6_v));
  assign n_829_v = ~(n_686_v);
  assign n_838_v = ~(n_2210_v);
  assign n_843_v = ~(n_2183_v);
  assign n_853_v = ~(v(n_525_v));
  assign n_855_v = ~((n_826_v|(n_844_v&n_2186_v)|(v(n_754_v)&(n_844_v|n_2186_v))));
  assign n_860_v = ~((n_811_v|v(n_856_v)));
  assign n_874_v = ~(n_877_v);
  assign n_877_v = ~((n_607_v|n_2278_v));
  assign n_882_v = ~(n_854_v);
  assign n_887_v = ~((v(n_892_v)|n_882_v|v(n_915_v)));
  assign n_888_v = ~(n_895_v);
  assign n_891_v = ~((v(n_892_v)|n_882_v));
  assign n_895_v = ~((n_2282_v|n_607_v));
  assign n_905_v = ~(v(n_2320_v));
  assign n_910_v = ~(n_911_v);
  assign n_911_v = ~((n_607_v|n_2394_v));
  assign n_926_v = ~(n_931_v);
  assign n_931_v = ~((n_2402_v|n_607_v));
  assign n_932_v = ~(n_842_v);
  assign n_939_v = ~(n_941_v);
  assign n_941_v = ~((n_607_v|n_2507_v));
  assign n_942_v = ~((v(n_950_v)|n_932_v|v(n_963_v)));
  assign n_955_v = ~((v(n_950_v)|v(n_963_v)|n_932_v|v(n_981_v)));
  assign n_961_v = ~(n_965_v);
  assign n_965_v = ~((n_2513_v|n_607_v));
  assign n_971_v = ~(v(n_2617_v));
  assign n_976_v = ~(n_977_v);
  assign n_977_v = ~((n_607_v|n_2614_v));
  assign n_987_v = ~(n_996_v);
  assign n_996_v = ~((n_2619_v|n_607_v));
  assign n_1012_v = ~(v(n_2700_v));
  assign n_1021_v = ~(v(n_2701_v));
  assign n_1022_v = ~(v(n_2702_v));
  assign n_1023_v = ~(v(n_2703_v));
  assign n_1024_v = ~(v(n_2704_v));
  assign n_1026_v = ~(v(n_1009_v));
  assign n_862_v = ~(n_762_v);
  assign n_866_v = ~(n_2227_v);
  assign n_869_v = ~(((n_2189_v&n_747_v)|(n_2226_v&n_831_v)));
  assign n_873_v = ~(v(n_755_v));
  assign n_875_v = ~((n_825_v|n_855_v));
  assign n_876_v = ~(v(n_861_v));
  assign n_890_v = ~(v(n_772_v));
  assign n_894_v = ~(n_2327_v);
  assign n_904_v = ~((n_826_v|(n_896_v&n_2330_v)|(n_878_v&(n_896_v|n_2330_v))));
  assign n_909_v = ~(v(n_783_v));
  assign n_919_v = ~(((n_2332_v&n_747_v)|(n_2390_v&n_831_v)));
  assign n_924_v = ~((n_825_v|n_904_v));
  assign n_927_v = ~(v(n_796_v));
  assign n_938_v = ~(v(n_803_v));
  assign n_940_v = ~(n_2493_v);
  assign n_952_v = ~((n_826_v|(n_943_v&n_2496_v)|(n_925_v&(n_943_v|n_2496_v))));
  assign n_962_v = ~(v(n_808_v));
  assign n_967_v = ~(((n_2498_v&n_747_v)|(n_2556_v&n_831_v)));
  assign n_972_v = ~((n_825_v|n_952_v));
  assign n_975_v = ~(v(n_836_v));
  assign n_986_v = ~(n_2657_v);
  assign n_990_v = ~(v(n_839_v));
  assign n_997_v = ~((n_826_v|(n_989_v&n_2659_v)|(n_767_v&(n_989_v|n_2659_v))));
  assign n_1006_v = ~(((n_2662_v&n_747_v)|(n_2682_v&n_831_v)));
  assign n_1008_v = ~((n_825_v|n_997_v));
  assign n_1010_v = ~(v(db4_v));
  assign n_1013_v = ~(v(n_1020_v));
  assign n_1015_v = ~(v(n_1014_v));
  assign n_1016_v = ~(v(n_1017_v));
  assign n_1019_v = ~(v(n_1018_v));
  assign n_1025_v = ~(v(n_2705_v));
  assign n_1047_v = ~(n_53_v);
  assign n_1046_v = ~((n_1041_v|v(clk_v)));
  assign n_1045_v = ~(n_63_v);
  assign n_1050_v = ~(n_83_v);
  assign n_1041_v = ~(n_1055_v);
  assign n_1057_v = ~((n_1052_v|n_63_v));
  assign n_1049_v = ~((v(clk_v)|n_102_v));
  assign n_1055_v = ~(n_1059_v);
  assign n_1065_v = ~(n_1057_v);
  assign n_1067_v = ~(v(_busrq_v));
  assign n_1071_v = ~(v(n_77_v));
  assign n_1086_v = ~(n_1067_v);
  assign n_1088_v = ~(n_64_v);
  assign n_1089_v = ~(v(_reset_v));
  assign n_1108_v = ~((v(n_81_v)|n_69_v));
  assign n_1091_v = ~((n_110_v|n_91_v));
  assign n_1093_v = ~(n_104_v);
  assign n_1094_v = ~(n_104_v);
  assign n_1097_v = ~(n_1089_v);
  assign n_1113_v = ~(v(n_128_v));
  assign n_1117_v = ~((n_69_v|v(n_120_v)));
  assign n_1125_v = ~(n_110_v);
  assign n_1106_v = ~(n_1105_v);
  assign n_1154_v = ~((n_105_v|v(n_92_v)));
  assign n_1132_v = ~((n_1124_v|n_103_v));
  assign n_1148_v = ~((n_1125_v|n_105_v));
  assign n_1137_v = ~((n_126_v|n_103_v|n_1146_v));
  assign n_1152_v = ~((n_126_v|n_1132_v));
  assign n_1151_v = ~((n_126_v|n_1133_v));
  assign n_1111_v = ~(n_1134_v);
  assign n_1146_v = ~(n_1135_v);
  assign n_1105_v = ~((n_1157_v&n_129_v));
  assign n_1144_v = ~(n_1137_v);
  assign n_1149_v = ~(n_1111_v);
  assign n_1123_v = ~(n_93_v);
  assign n_1156_v = ~(n_1155_v);
  assign n_1165_v = ~((n_141_v&n_54_v));
  assign n_1153_v = ~((n_1159_v&n_129_v));
  assign n_1141_v = ~((n_1174_v|v(clk_v)));
  assign n_1187_v = ~((_t3_v|n_95_v));
  assign n_1173_v = ~((v(n_127_v)|_t2_v));
  assign n_1143_v = ~(n_1153_v);
  assign n_1191_v = ~(v(n_89_v));
  assign n_1177_v = ~((n_1183_v&n_129_v));
  assign n_1179_v = ~(n_1152_v);
  assign n_1133_v = ~(n_1192_v);
  assign n_1194_v = ~(v(n_1170_v));
  assign n_1155_v = ~((n_72_v|v(n_157_v)));
  assign n_1186_v = ~(n_184_v);
  assign n_1197_v = ~(v(n_147_v));
  assign n_1190_v = ~(n_1201_v);
  assign n_1205_v = ~((m1_v&_t2_v));
  assign n_1209_v = ~(v(n_140_v));
  assign n_1201_v = ~((n_1212_v&n_129_v));
  assign n_1216_v = ~((v(n_176_v)|v(n_118_v)));
  assign n_1208_v = ~(((m1_v&_t2_v)|(_t1_v&(n_193_v&m3_v))));
  assign n_1213_v = ~(n_1238_v);
  assign n_1236_v = ~(v(n_1228_v));
  assign n_1241_v = ~(v(n_1225_v));
  assign n_1238_v = ~((n_126_v|n_1250_v|n_103_v));
  assign n_1252_v = ~((m1_v&_t2_v));
  assign n_1249_v = ~(v(n_185_v));
  assign n_1247_v = ~(v(n_1221_v));
  assign n_1250_v = ~(n_1258_v);
  assign n_1266_v = ~(n_1261_v);
  assign n_1286_v = ~((n_1251_v|v(clk_v)));
  assign n_1256_v = ~(n_192_v);
  assign n_1233_v = ~(n_198_v);
  assign n_1276_v = ~(((_t2_v|v(n_223_v))&(n_177_v|(m1_v&n_188_v))));
  assign n_1281_v = ~((n_212_v&(m2_v|(n_202_v&m1_v))));
  assign n_1270_v = ~(n_1272_v);
  assign n_1265_v = ~((n_1266_v|v(clk_v)));
  assign n_1292_v = ~((n_95_v|n_215_v));
  assign n_1295_v = ~(v(n_1271_v));
  assign n_1294_v = ~(n_308_v);
  assign n_1293_v = ~(n_224_v);
  assign n_1304_v = ~(n_238_v);
  assign n_1298_v = ~((n_234_v|n_213_v));
  assign n_1314_v = ~(n_208_v);
  assign n_1318_v = ~(n_252_v);
  assign n_1322_v = ~(n_110_v);
  assign n_1315_v = ~(n_246_v);
  assign n_1326_v = ~(n_1323_v);
  assign n_1328_v = ~(n_1334_v);
  assign n_1333_v = ~(n_211_v);
  assign n_1335_v = ~((v(clk_v)|n_1326_v));
  assign n_1285_v = ~((v(n_190_v)|n_1337_v));
  assign n_1334_v = ~(n_1342_v);
  assign n_1339_v = ~(v(n_240_v));
  assign n_1337_v = ~(n_239_v);
  assign n_1345_v = ~((n_95_v|_t1_v));
  assign n_1344_v = ~(v(n_259_v));
  assign n_1346_v = ~(v(n_216_v));
  assign n_1351_v = ~(n_260_v);
  assign n_1353_v = ~(n_110_v);
  assign n_1352_v = ~(n_360_v);
  assign n_1357_v = ~(n_1356_v);
  assign n_1355_v = ~(n_318_v);
  assign n_1361_v = ~((m4_v|(n_329_v&m3_v)));
  assign n_1381_v = ~((n_65_v|n_390_v));
  assign n_1382_v = ~(n_194_v);
  assign n_1389_v = ~((n_391_v|(n_395_v&n_1382_v)));
  assign n_1392_v = ~(n_396_v);
  assign n_1391_v = ~(n_1384_v);
  assign n_1384_v = ~(n_1398_v);
  assign n_1397_v = ~((n_262_v|n_330_v));
  assign n_1396_v = ~(n_1397_v);
  assign n_1399_v = ~((n_401_v|n_416_v));
  assign n_1401_v = ~(n_371_v);
  assign n_1402_v = ~(n_381_v);
  assign n_1403_v = ~(n_420_v);
  assign n_1406_v = ~((n_419_v|n_385_v));
  assign n_1410_v = ~(n_1404_v);
  assign n_1413_v = ~((n_407_v&n_1411_v));
  assign n_1411_v = ~((_t1_v&((n_1406_v&m3_v)|(m4_v&(n_387_v&n_395_v))|(m2_v&(n_1406_v|n_270_v)))));
  assign n_1404_v = ~(n_1414_v);
  assign n_1415_v = ~((n_419_v&(n_232_v|n_220_v)));
  assign n_1412_v = ~((n_228_v|n_270_v));
  assign n_1418_v = ~(v(n_408_v));
  assign n_1420_v = ~(((_t2_v&((n_1415_v&m4_v)|(n_1417_v&m2_v)))|(_t4_v&(m5_v|((n_262_v|n_395_v)&(m4_v|m3_v))))));
  assign n_1421_v = ~(n_467_v);
  assign n_1417_v = ~((n_419_v&n_1425_v));
  assign n_1432_v = ~((n_1420_v&n_440_v));
  assign n_1427_v = ~((n_95_v|(n_1426_v&(m1_v&_t1_v))));
  assign n_1430_v = ~(n_327_v);
  assign n_1431_v = ~(n_1427_v);
  assign n_1425_v = ~((n_270_v|n_318_v));
  assign n_1426_v = ~(n_99_v);
  assign n_1442_v = ~(n_1433_v);
  assign n_1434_v = ~(n_387_v);
  assign n_1448_v = ~(n_232_v);
  assign n_1465_v = ~((n_232_v|n_417_v));
  assign n_1444_v = ~((n_361_v|n_261_v));
  assign n_1463_v = ~(n_417_v);
  assign n_1458_v = ~((n_459_v|n_398_v));
  assign n_1445_v = ~((n_488_v|n_446_v));
  assign n_1450_v = ~(n_1445_v);
  assign n_1455_v = ~(n_424_v);
  assign n_1451_v = ~(n_1442_v);
  assign n_1474_v = ~((n_192_v|n_232_v));
  assign n_1449_v = ~(n_453_v);
  assign n_1464_v = ~(n_202_v);
  assign n_1471_v = ~(n_1440_v);
  assign n_1476_v = ~(n_110_v);
  assign n_1479_v = ~((n_1432_v|n_465_v));
  assign n_1477_v = ~((n_466_v|n_1464_v));
  assign n_1475_v = ~((n_467_v|n_1478_v));
  assign n_1490_v = ~(n_441_v);
  assign n_1489_v = ~(n_435_v);
  assign n_1484_v = ~((n_478_v|n_464_v));
  assign n_1480_v = ~(n_262_v);
  assign n_1481_v = ~(n_461_v);
  assign n_1478_v = ~(n_456_v);
  assign n_1504_v = ~(n_1499_v);
  assign n_1500_v = ~(n_1484_v);
  assign n_1503_v = ~((n_1480_v|n_324_v));
  assign n_1502_v = ~(n_220_v);
  assign n_1505_v = ~(n_1504_v);
  assign n_1509_v = ~(n_101_v);
  assign n_1506_v = ~(n_270_v);
  assign n_1508_v = ~((n_398_v|n_194_v));
  assign n_1511_v = ~(n_493_v);
  assign n_1513_v = ~(n_1512_v);
  assign n_1514_v = ~(n_1513_v);
  assign n_1522_v = ~(n_473_v);
  assign n_1533_v = ~(n_514_v);
  assign n_1541_v = ~(((_t3_v&(n_1475_v&(m5_v|m4_v)))|((n_318_v|n_446_v|n_330_v)&(_t1_v&(m5_v|m4_v)))));
  assign n_1553_v = ~((n_320_v&((m2_v&_t3_v)|(m3_v&_t2_v))));
  assign n_1561_v = ~((((n_270_v|n_434_v)&(m3_v&_t2_v))|(_t3_v&((n_492_v&m4_v)|(m2_v&(n_1450_v&n_1506_v))))));
  assign n_1556_v = ~(((_t4_v&(n_315_v&m1_v))|(_t3_v&(n_270_v&m2_v))));
  assign n_1552_v = ~((((n_395_v|n_334_v)&(m1_v&_t5_v))|(_t2_v&((n_395_v&(m3_v|m4_v))|(m5_v&(n_456_v&n_395_v))))));
  assign n_1554_v = ~(((_t1_v&(n_1500_v&m2_v))|(_t3_v&((n_492_v&m5_v)|(n_1450_v&m3_v)))));
  assign n_1557_v = ~(((_t3_v|_t1_v)&(n_289_v&(m5_v|m4_v))));
  assign n_1550_v = ~((m1_v&_t2_v));
  assign n_1592_v = ~(n_1575_v);
  assign n_1551_v = ~((n_333_v&n_535_v));
  assign n_1573_v = ~((n_1553_v&(n_555_v|n_1601_v|n_484_v)));
  assign n_1576_v = ~(n_1557_v);
  assign n_1582_v = ~((n_504_v&(n_555_v&n_529_v)));
  assign n_1593_v = ~(n_1602_v);
  assign n_1583_v = ~(n_1474_v);
  assign n_1584_v = ~(n_508_v);
  assign n_1578_v = ~((n_507_v&n_506_v));
  assign n_1580_v = ~(n_1553_v);
  assign n_1607_v = ~(n_1592_v);
  assign n_1577_v = ~((n_1597_v|n_578_v));
  assign n_1585_v = ~((n_512_v&n_1554_v));
  assign n_1599_v = ~(n_520_v);
  assign n_1609_v = ~(n_66_v);
  assign n_1645_v = ~(n_559_v);
  assign n_1629_v = ~((n_479_v|n_568_v));
  assign n_1605_v = ~(n_505_v);
  assign n_1643_v = ~((n_548_v|n_484_v));
  assign n_1641_v = ~((n_1585_v|(n_585_v&(n_479_v|n_568_v))));
  assign n_1628_v = ~((n_1550_v&n_547_v));
  assign n_1646_v = ~((n_548_v|n_563_v));
  assign n_1608_v = ~(n_484_v);
  assign n_1621_v = ~((n_1556_v&(n_547_v&n_1550_v)));
  assign n_1635_v = ~(n_1577_v);
  assign n_1648_v = ~((n_1621_v|n_95_v));
  assign n_1636_v = ~(n_555_v);
  assign n_1601_v = ~(n_548_v);
  assign n_1616_v = ~((n_518_v&n_567_v));
  assign n_1640_v = ~(n_1655_v);
  assign n_1644_v = ~(n_1630_v);
  assign n_1647_v = ~((n_532_v|(n_1629_v&n_585_v)|(n_571_v&n_558_v)));
  assign n_1651_v = ~(n_1650_v);
  assign n_1650_v = ~(n_580_v);
  assign n_1632_v = ~((v(n_562_v)|(n_1609_v&v(clk_v))));
  assign n_1656_v = ~(n_1667_v);
  assign n_1665_v = ~((v(n_562_v)|(n_1609_v&v(clk_v))));
  assign n_1655_v = ~(n_1615_v);
  assign n_1657_v = ~(n_1663_v);
  assign n_1658_v = ~(n_578_v);
  assign n_1703_v = ~(n_1675_v);
  assign n_1687_v = ~(n_1676_v);
  assign n_1716_v = ~((v(clk_v)|n_519_v));
  assign n_1707_v = ~(n_1685_v);
  assign n_1713_v = ~(ex_dehl_combined_v);
  assign n_1708_v = ~(ex_dehl_combined_v);
  assign n_1711_v = ~(n_591_v);
  assign n_1712_v = ~(n_1705_v);
  assign n_1714_v = ~(n_1706_v);
  assign n_1715_v = ~(n_1656_v);
  assign n_1717_v = ~(n_1695_v);
  assign n_1737_v = ~(n_393_v);
  assign n_1725_v = ~(n_1733_v);
  assign n_1736_v = ~((n_685_v|n_651_v));
  assign n_1733_v = ~(v(clk_v));
  assign n_1695_v = ~(n_1725_v);
  assign n_1738_v = ~((n_1711_v&n_630_v));
  assign n_1739_v = ~((n_591_v&n_630_v));
  assign n_1740_v = ~((n_640_v&n_1712_v));
  assign n_1741_v = ~((n_634_v&n_1712_v));
  assign n_1742_v = ~((n_640_v&n_1714_v));
  assign n_1743_v = ~((n_634_v&n_1714_v));
  assign n_1744_v = ~((n_640_v&n_1715_v));
  assign n_1745_v = ~((n_634_v&n_1715_v));
  assign n_1746_v = ~((v(n_633_v)&n_1657_v));
  assign n_1747_v = ~((n_1657_v&v(ex_af_v)));
  assign n_1722_v = ~((n_534_v|n_634_v|v(clk_v)));
  assign n_1719_v = ~((n_640_v|n_534_v|v(clk_v)));
  assign n_1779_v = ~((n_1774_v|n_627_v));
  assign n_1777_v = ~(n_1776_v);
  assign n_1795_v = ~((n_588_v|v(clk_v)));
  assign n_1796_v = ~((n_590_v|v(clk_v)));
  assign n_1797_v = ~((n_1674_v|v(clk_v)));
  assign n_1803_v = ~((n_589_v|v(clk_v)));
  assign n_1804_v = ~((v(n_689_v)|n_627_v));
  assign n_1774_v = ~(v(n_689_v));
  assign n_1828_v = ~(v(n_703_v));
  assign n_1776_v = ~(n_1830_v);
  assign n_1835_v = ~(n_1776_v);
  assign n_1832_v = ~(n_1776_v);
  assign n_1829_v = ~(n_1774_v);
  assign n_1834_v = ~(n_1776_v);
  assign n_1836_v = ~((n_406_v|v(n_709_v)));
  assign n_1856_v = ~(n_1776_v);
  assign n_1840_v = ~(n_436_v);
  assign n_1837_v = ~(n_694_v);
  assign n_1884_v = ~((n_627_v|v(n_723_v)));
  assign n_1865_v = ~(n_436_v);
  assign n_1866_v = ~(n_1836_v);
  assign n_1887_v = ~(n_1886_v);
  assign n_1889_v = ~(n_1886_v);
  assign n_1907_v = ~(n_1910_v);
  assign n_1888_v = ~(n_1886_v);
  assign n_1886_v = ~(n_1909_v);
  assign n_1883_v = ~(n_1886_v);
  assign n_1906_v = ~(v(n_731_v));
  assign n_1929_v = ~(v(n_739_v));
  assign n_1914_v = ~(n_1931_v);
  assign n_1910_v = ~(v(n_723_v));
  assign n_1937_v = ~(n_1914_v);
  assign n_1934_v = ~(n_1914_v);
  assign n_1936_v = ~(n_1914_v);
  assign n_1938_v = ~((n_730_v|v(n_746_v)));
  assign n_1941_v = ~(n_436_v);
  assign n_1963_v = ~(n_1914_v);
  assign n_1939_v = ~(n_710_v);
  assign n_1971_v = ~(n_1938_v);
  assign n_1988_v = ~(n_436_v);
  assign n_1969_v = ~((n_1910_v|n_627_v));
  assign n_1993_v = ~(n_1992_v);
  assign n_1995_v = ~(n_1992_v);
  assign n_1994_v = ~(n_1992_v);
  assign n_1992_v = ~(n_2013_v);
  assign n_1990_v = ~(n_1992_v);
  assign n_2012_v = ~(v(n_774_v));
  assign n_2014_v = ~((n_627_v|n_778_v));
  assign n_2033_v = ~(v(n_777_v));
  assign n_2018_v = ~(n_2034_v);
  assign n_2038_v = ~(n_2018_v);
  assign n_2035_v = ~(n_2018_v);
  assign n_2037_v = ~(n_2018_v);
  assign n_2039_v = ~((n_773_v|v(n_787_v)));
  assign n_2042_v = ~(n_436_v);
  assign n_2060_v = ~(n_2018_v);
  assign n_2040_v = ~(n_748_v);
  assign n_2067_v = ~(n_2039_v);
  assign n_2085_v = ~(n_436_v);
  assign n_2089_v = ~(n_2088_v);
  assign n_2093_v = ~(n_2088_v);
  assign n_2092_v = ~(n_2088_v);
  assign n_2088_v = ~(n_2114_v);
  assign n_2086_v = ~(n_2088_v);
  assign n_2113_v = ~(v(n_806_v));
  assign n_2133_v = ~(v(n_810_v));
  assign n_2118_v = ~(n_2134_v);
  assign n_2138_v = ~(n_2118_v);
  assign n_2135_v = ~(n_2118_v);
  assign n_2137_v = ~(n_2118_v);
  assign n_2117_v = ~((v(n_2116_v)|n_627_v));
  assign n_2141_v = ~(n_436_v);
  assign n_2157_v = ~(n_2118_v);
  assign n_2139_v = ~(n_789_v);
  assign n_2164_v = ~(n_690_v);
  assign n_2180_v = ~(n_436_v);
  assign n_2190_v = ~(n_2187_v);
  assign n_2220_v = ~(n_778_v);
  assign n_2195_v = ~(n_2187_v);
  assign n_2194_v = ~(n_2187_v);
  assign n_2187_v = ~(n_2222_v);
  assign n_2182_v = ~(n_2187_v);
  assign n_2221_v = ~(v(n_863_v));
  assign n_2246_v = ~(v(n_871_v));
  assign n_2225_v = ~(n_2248_v);
  assign n_2252_v = ~(n_2225_v);
  assign n_2249_v = ~(n_2225_v);
  assign n_2251_v = ~(n_2225_v);
  assign n_2257_v = ~(n_436_v);
  assign n_2275_v = ~(n_2225_v);
  assign n_2253_v = ~(n_860_v);
  assign n_2281_v = ~(n_854_v);
  assign n_2298_v = ~(n_436_v);
  assign n_2303_v = ~(n_2301_v);
  assign n_2302_v = ~(n_905_v);
  assign n_2305_v = ~(n_2301_v);
  assign n_2304_v = ~(n_2301_v);
  assign n_2301_v = ~(n_2329_v);
  assign n_2299_v = ~(n_2301_v);
  assign n_2325_v = ~(v(n_901_v));
  assign n_2359_v = ~(v(n_907_v));
  assign n_2343_v = ~(n_2361_v);
  assign n_2365_v = ~(n_2343_v);
  assign n_2362_v = ~(n_2343_v);
  assign n_2364_v = ~(n_2343_v);
  assign n_2386_v = ~((n_627_v|v(n_2320_v)));
  assign n_2368_v = ~(n_436_v);
  assign n_2387_v = ~(n_2343_v);
  assign n_2366_v = ~(n_891_v);
  assign n_2401_v = ~(n_887_v);
  assign n_2418_v = ~(n_436_v);
  assign n_2424_v = ~(n_2422_v);
  assign n_2428_v = ~(n_2422_v);
  assign n_2427_v = ~(n_2422_v);
  assign n_2422_v = ~(n_2448_v);
  assign n_2419_v = ~(n_2422_v);
  assign n_2446_v = ~(v(n_933_v));
  assign n_2464_v = ~(v(n_936_v));
  assign n_2449_v = ~(n_2465_v);
  assign n_2469_v = ~(n_2449_v);
  assign n_2466_v = ~(n_2449_v);
  assign n_2468_v = ~(n_2449_v);
  assign n_2472_v = ~((v(n_950_v)|n_932_v));
  assign n_2473_v = ~(n_436_v);
  assign n_2495_v = ~(n_2449_v);
  assign n_2470_v = ~(n_842_v);
  assign n_2506_v = ~((n_905_v|n_627_v));
  assign n_2512_v = ~(n_2472_v);
  assign n_2529_v = ~(n_436_v);
  assign n_2536_v = ~(n_2534_v);
  assign n_2553_v = ~((n_627_v|n_971_v));
  assign n_2538_v = ~(n_2534_v);
  assign n_2537_v = ~(n_2534_v);
  assign n_2534_v = ~(n_2562_v);
  assign n_2532_v = ~(n_2534_v);
  assign n_2559_v = ~(v(n_969_v));
  assign n_2587_v = ~(v(n_974_v));
  assign n_2572_v = ~(n_2588_v);
  assign n_2592_v = ~(n_2572_v);
  assign n_2589_v = ~(n_2572_v);
  assign n_2591_v = ~(n_2572_v);
  assign n_2596_v = ~(n_436_v);
  assign n_2612_v = ~(n_2572_v);
  assign n_2593_v = ~(n_942_v);
  assign n_2618_v = ~(n_955_v);
  assign n_2640_v = ~(n_2660_v);
  assign n_2636_v = ~((v(n_2617_v)|n_627_v));
  assign n_2642_v = ~(n_2660_v);
  assign n_2639_v = ~(n_2660_v);
  assign n_2660_v = ~(n_2674_v);
  assign n_2671_v = ~(v(n_998_v));
  assign n_2689_v = ~(n_971_v);
  assign n_2698_v = ~(n_1026_v);
  assign n_2696_v = ~((v(n_1009_v)|n_627_v));
  assign n_2708_v = ~((n_627_v|n_1026_v));
  assign n_2725_v = ~((v(n_2700_v)|n_627_v));
  assign n_2719_v = ~((n_1012_v|n_627_v));
  assign n_2727_v = ~((n_627_v|v(n_2701_v)));
  assign n_2728_v = ~((v(n_2702_v)|n_627_v));
  assign n_2729_v = ~((n_627_v|v(n_2703_v)));
  assign n_2730_v = ~((v(n_2704_v)|n_627_v));
  assign n_2710_v = ~((n_627_v|n_1021_v));
  assign n_2711_v = ~((n_627_v|n_1022_v));
  assign n_2712_v = ~((n_627_v|n_1023_v));
  assign n_2713_v = ~((n_627_v|n_1024_v));
  assign n_2715_v = ~(n_1012_v);
  assign n_2720_v = ~(n_1021_v);
  assign n_2721_v = ~(n_1022_v);
  assign n_2722_v = ~(n_1023_v);
  assign n_2723_v = ~(n_1024_v);
  assign n_1056_v = ~((n_60_v|n_1048_v));
  assign n_1054_v = ~(n_60_v);
  assign n_1048_v = ~(n_1054_v);
  assign n_1066_v = ~(n_80_v);
  assign n_1064_v = ~(v(n_84_v));
  assign n_1063_v = ~(n_108_v);
  assign n_1073_v = ~(v(_int_v));
  assign n_1069_v = ~(v(n_1072_v));
  assign n_1074_v = ~((n_69_v|v(n_85_v)));
  assign n_1075_v = ~(v(n_1077_v));
  assign n_1068_v = ~(n_1073_v);
  assign n_1070_v = ~((n_113_v|(n_79_v&n_122_v)));
  assign n_1085_v = ~((n_154_v&(n_188_v&m1_v)));
  assign n_1104_v = ~((n_69_v|v(n_86_v)));
  assign n_1103_v = ~(v(n_1076_v));
  assign n_1083_v = ~((n_1096_v|v(clk_v)));
  assign n_1100_v = ~((n_1107_v|n_188_v));
  assign n_1087_v = ~((n_1109_v|n_109_v));
  assign n_1110_v = ~(n_114_v);
  assign n_1116_v = ~(n_79_v);
  assign n_1112_v = ~(n_99_v);
  assign n_1115_v = ~(n_101_v);
  assign n_1120_v = ~((n_121_v|v(clk_v)));
  assign n_1119_v = ~(n_1140_v);
  assign n_1139_v = ~((n_107_v&_t1_v));
  assign n_1131_v = ~(((_t1_v&n_1142_v)|(m1_v&(_t3_v|(_t1_v&n_1164_v)))));
  assign n_1130_v = ~((n_1147_v|v(clk_v)));
  assign n_1128_v = ~((n_1158_v|v(clk_v)));
  assign n_1127_v = ~(n_106_v);
  assign n_1150_v = ~(v(db0_v));
  assign n_1118_v = ~(v(n_1126_v));
  assign n_1081_v = ~((v(clk_v)|n_1160_v));
  assign n_1109_v = ~(n_1163_v);
  assign n_1166_v = ~(n_231_v);
  assign n_1182_v = ~(n_1167_v);
  assign n_1167_v = ~(n_1145_v);
  assign n_1172_v = ~(n_1162_v);
  assign n_1082_v = ~(n_1169_v);
  assign n_1121_v = ~((n_1175_v|n_1176_v));
  assign n_1140_v = ~((v(clk_v)&(m1_v&_t3_v)));
  assign n_1169_v = ~((_t3_v&m1_v));
  assign n_1175_v = ~(n_177_v);
  assign n_1195_v = ~((n_156_v&n_1172_v));
  assign n_1188_v = ~(n_142_v);
  assign n_1189_v = ~((n_142_v&(n_188_v&n_1180_v)));
  assign n_1198_v = ~((_t2_v&n_177_v));
  assign n_1193_v = ~(v(n_149_v));
  assign n_1181_v = ~(n_117_v);
  assign n_1176_v = ~((_t2_v&n_107_v));
  assign n_1199_v = ~((n_95_v|(n_1229_v&_t3_v)));
  assign n_1196_v = ~((n_133_v|n_82_v));
  assign n_1202_v = ~((n_1195_v|v(clk_v)));
  assign n_1203_v = ~((n_165_v|n_123_v));
  assign n_1136_v = ~(n_236_v);
  assign n_1084_v = ~(n_1198_v);
  assign n_1185_v = ~(_t2_v);
  assign n_1206_v = ~((_t1_v&(n_249_v&m1_v)));
  assign n_1211_v = ~(n_179_v);
  assign n_1246_v = ~(((_t4_v|n_95_v)|(_t3_v&n_1231_v)));
  assign n_1214_v = ~((n_178_v|n_204_v));
  assign n_1210_v = ~(n_191_v);
  assign n_1164_v = ~(n_188_v);
  assign n_1215_v = ~(n_1211_v);
  assign n_1142_v = ~((n_177_v|m1_v));
  assign n_1099_v = ~(n_258_v);
  assign n_1180_v = ~((n_236_v|n_218_v));
  assign n_1226_v = ~((n_170_v|n_165_v));
  assign n_1147_v = ~(n_1235_v);
  assign n_1223_v = ~(v(n_1220_v));
  assign n_1224_v = ~((_t2_v&(n_237_v&m1_v)));
  assign n_1239_v = ~(n_1278_v);
  assign n_1255_v = ~((n_1243_v|(n_200_v&n_204_v)));
  assign n_1248_v = ~(n_1331_v);
  assign n_1262_v = ~(n_1254_v);
  assign n_1259_v = ~(n_1245_v);
  assign n_1254_v = ~(n_1242_v);
  assign n_1267_v = ~(n_1255_v);
  assign n_1257_v = ~(v(db1_v));
  assign n_1273_v = ~(n_1259_v);
  assign n_1274_v = ~(n_1246_v);
  assign n_1282_v = ~(((_t1_v&n_107_v)|(_t3_v&(n_1263_v&n_125_v))));
  assign n_1231_v = ~(m1_v);
  assign n_1260_v = ~((n_142_v&(n_188_v&n_218_v)));
  assign n_1280_v = ~(n_182_v);
  assign n_1275_v = ~((_t2_v&m1_v));
  assign n_1278_v = ~(n_206_v);
  assign n_1297_v = ~((n_1267_v|n_204_v));
  assign n_1287_v = ~((n_188_v&n_218_v));
  assign n_1277_v = ~(n_205_v);
  assign n_1283_v = ~((_t1_v&(m1_v&n_245_v)));
  assign n_1229_v = ~(m1_v);
  assign n_1284_v = ~((n_135_v&n_142_v));
  assign n_1299_v = ~((n_1167_v|n_1279_v));
  assign n_1268_v = ~(n_1277_v);
  assign n_1291_v = ~((n_95_v|_t3_v));
  assign n_1279_v = ~(n_201_v);
  assign n_1289_v = ~(n_1189_v);
  assign n_1263_v = ~((m1_v|(n_164_v&m3_v)|(m3_v&n_193_v)));
  assign n_1296_v = ~(n_1319_v);
  assign n_1290_v = ~(n_195_v);
  assign n_1301_v = ~(n_1282_v);
  assign n_1288_v = ~(n_1290_v);
  assign n_1303_v = ~(n_1259_v);
  assign n_1264_v = ~(n_1310_v);
  assign n_1311_v = ~((m3_v&(_t3_v&n_193_v)));
  assign n_1308_v = ~((n_133_v|n_82_v));
  assign n_1312_v = ~(n_1254_v);
  assign n_1309_v = ~(n_226_v);
  assign n_1310_v = ~(n_1321_v);
  assign n_1237_v = ~((n_1287_v|n_236_v));
  assign n_1317_v = ~(n_1299_v);
  assign n_1305_v = ~(n_228_v);
  assign n_1316_v = ~(n_1297_v);
  assign n_1330_v = ~((n_165_v|n_195_v));
  assign n_1325_v = ~((n_311_v|n_312_v));
  assign n_1340_v = ~((n_255_v|v(n_244_v)));
  assign n_1338_v = ~((n_165_v|n_250_v));
  assign n_1349_v = ~(v(db7_v));
  assign n_1348_v = ~(n_1350_v);
  assign n_1359_v = ~(n_1360_v);
  assign n_1363_v = ~(n_358_v);
  assign n_1365_v = ~(n_1366_v);
  assign n_1362_v = ~(n_1363_v);
  assign n_1369_v = ~(n_1370_v);
  assign n_1367_v = ~((n_133_v|n_82_v));
  assign n_1372_v = ~((n_165_v|n_358_v));
  assign n_1374_v = ~(n_1375_v);
  assign n_1378_v = ~((n_165_v|n_383_v));
  assign n_1379_v = ~(n_1380_v);
  assign n_1387_v = ~(n_1388_v);
  assign n_1394_v = ~(n_1395_v);
  assign n_1400_v = ~(n_326_v);
  assign n_1407_v = ~((n_133_v|n_82_v));
  assign n_1408_v = ~(n_1409_v);
  assign n_1409_v = ~(n_414_v);
  assign n_1419_v = ~(n_1416_v);
  assign n_1424_v = ~(n_348_v);
  assign n_1423_v = ~(n_1419_v);
  assign n_1422_v = ~(v(db2_v));
  assign n_1429_v = ~((n_344_v|n_299_v));
  assign n_1428_v = ~((n_165_v|n_414_v));
  assign n_1456_v = ~(n_403_v);
  assign n_1441_v = ~((n_165_v|n_452_v));
  assign n_1446_v = ~(n_247_v);
  assign n_1467_v = ~((n_272_v|n_349_v));
  assign n_1454_v = ~((n_273_v|n_350_v));
  assign n_1459_v = ~(n_423_v);
  assign n_1453_v = ~((n_330_v|n_446_v));
  assign n_1472_v = ~(((n_378_v&n_450_v)|(n_1393_v&n_447_v)));
  assign n_1468_v = ~(((n_375_v&n_450_v)|(n_1446_v&n_447_v)));
  assign n_1469_v = ~(((n_374_v&n_450_v)|(n_449_v&n_447_v)));
  assign n_1443_v = ~((n_272_v&n_449_v));
  assign n_1461_v = ~(n_421_v);
  assign n_1457_v = ~(n_409_v);
  assign n_1447_v = ~(n_428_v);
  assign n_1452_v = ~((n_469_v&n_254_v));
  assign n_1460_v = ~(n_1438_v);
  assign n_1470_v = ~(((n_330_v|n_228_v)|(n_488_v&n_456_v)));
  assign n_1473_v = ~(n_425_v);
  assign n_1486_v = ~(n_415_v);
  assign n_1493_v = ~(n_1452_v);
  assign n_1494_v = ~(n_405_v);
  assign n_1487_v = ~(n_270_v);
  assign n_1483_v = ~(n_444_v);
  assign n_1485_v = ~(n_404_v);
  assign n_1482_v = ~(n_1469_v);
  assign n_1488_v = ~(n_1429_v);
  assign n_1492_v = ~(n_1472_v);
  assign n_1495_v = ~(n_1468_v);
  assign n_1496_v = ~(n_352_v);
  assign n_1497_v = ~(n_1467_v);
  assign n_1510_v = ~((n_87_v|n_487_v));
  assign n_1518_v = ~((_t3_v&(n_220_v&m2_v)));
  assign n_1516_v = ~((n_222_v|(n_1515_v&(m1_v&_t5_v))));
  assign n_1517_v = ~((n_1456_v&((m4_v&_t3_v)|(m1_v&_t4_v))));
  assign n_1520_v = ~(((_t1_v&(n_271_v&m4_v))|(_t3_v&((n_228_v&m4_v)|(m3_v&(n_271_v|n_270_v))))));
  assign n_1521_v = ~(((m1_v&_t4_v)|((n_469_v|n_463_v)&(m4_v&_t3_v))));
  assign n_1519_v = ~((((_t5_v&(n_228_v&m1_v))|(_t3_v&(m1_v|m2_v)))|(_t1_v&((n_330_v&m5_v)|(m4_v&(n_330_v|n_469_v))))));
  assign n_1532_v = ~(((m1_v&_t3_v)|((n_469_v|n_463_v)&(m4_v&_t2_v))));
  assign n_1526_v = ~((((m1_v&_t5_v)|(_t2_v&(n_330_v&m5_v)))|(_t1_v&((n_439_v&m1_v)|(m3_v&(n_323_v|n_220_v))))));
  assign n_1525_v = ~(((_t1_v&(n_1493_v&m4_v))|(_t3_v&(n_254_v&m1_v))));
  assign n_1524_v = ~((_t5_v&(n_229_v&m1_v)));
  assign n_1529_v = ~(((m1_v&_t4_v)|(m2_v&_t2_v)|(m4_v&_t1_v)));
  assign n_1534_v = ~(((_t4_v&(n_366_v&m1_v))|(_t1_v&(n_1487_v&m3_v))));
  assign n_1530_v = ~((_t1_v&(m1_v&(n_470_v|n_1485_v))));
  assign n_1515_v = ~(((n_352_v|n_219_v)&(_t4_v|_t5_v)));
  assign n_1523_v = ~((_t2_v&(n_1457_v&m1_v)));
  assign n_1531_v = ~((_t3_v&(n_220_v&m2_v)));
  assign n_1528_v = ~(((n_353_v&m2_v)|(m3_v&(n_322_v|n_323_v))));
  assign n_1538_v = ~(n_1521_v);
  assign n_1539_v = ~(n_1525_v);
  assign n_1540_v = ~(n_1520_v);
  assign n_1546_v = ~((_t1_v&(n_296_v&m1_v)));
  assign n_1542_v = ~((n_1524_v&n_496_v));
  assign n_1558_v = ~(((_t3_v&(n_220_v&m3_v))|(_t1_v&((n_491_v&m5_v)|(m4_v&(n_488_v|n_478_v))))));
  assign n_1536_v = ~(n_1527_v);
  assign n_1544_v = ~((n_524_v&n_463_v));
  assign n_1545_v = ~(n_1524_v);
  assign n_1574_v = ~(n_460_v);
  assign n_1572_v = ~((n_1543_v|n_1549_v));
  assign n_1548_v = ~(n_503_v);
  assign n_1571_v = ~(n_1534_v);
  assign n_1594_v = ~(n_1547_v);
  assign n_1591_v = ~((n_1555_v|v(clk_v)));
  assign n_1588_v = ~(n_1516_v);
  assign n_1595_v = ~((n_1559_v|n_1540_v));
  assign n_1579_v = ~((n_543_v|v(clk_v)));
  assign n_1581_v = ~(n_1535_v);
  assign n_1596_v = ~(n_498_v);
  assign n_1587_v = ~(n_1568_v);
  assign n_1598_v = ~(n_1567_v);
  assign n_1606_v = ~(n_1570_v);
  assign n_1566_v = ~(n_515_v);
  assign n_1600_v = ~(n_1569_v);
  assign n_1589_v = ~((n_533_v&n_523_v));
  assign n_1565_v = ~((n_1610_v&n_550_v));
  assign n_1633_v = ~((n_1589_v|(n_554_v&n_556_v)|(n_549_v&n_558_v)));
  assign n_1623_v = ~(n_1515_v);
  assign n_1617_v = ~(n_1603_v);
  assign n_1624_v = ~(n_530_v);
  assign n_1622_v = ~(n_306_v);
  assign n_1618_v = ~(n_1523_v);
  assign n_1619_v = ~((n_1612_v|n_1581_v));
  assign n_1625_v = ~(n_1587_v);
  assign n_1627_v = ~(n_1532_v);
  assign n_1634_v = ~(n_1565_v);
  assign n_1620_v = ~(n_1595_v);
  assign n_1642_v = ~(n_1606_v);
  assign n_1626_v = ~(v(n_1586_v));
  assign n_1638_v = ~(n_1598_v);
  assign n_1631_v = ~(n_1600_v);
  assign n_1639_v = ~(n_1637_v);
  assign n_1662_v = ~((n_1624_v|n_561_v));
  assign n_1654_v = ~((n_1652_v&n_582_v));
  assign n_1612_v = ~(n_1660_v);
  assign n_1668_v = ~((n_583_v|n_1659_v));
  assign n_1661_v = ~(n_598_v);
  assign n_1680_v = ~((n_1654_v|v(clk_v)));
  assign n_1686_v = ~(((m3_v&_t3_v)|(_t4_v&(n_330_v&m4_v))));
  assign n_1637_v = ~(n_1673_v);
  assign n_1698_v = ~((m3_v&(_t5_v|_t4_v|_t3_v)));
  assign n_1690_v = ~(((_t2_v&(n_330_v&m4_v))|(_t4_v&(n_220_v&(m4_v|m3_v)))));
  assign n_1671_v = ~(n_558_v);
  assign n_1684_v = ~((_t4_v|_t2_v));
  assign n_1689_v = ~(((_t2_v&(n_220_v&m3_v))|(_t3_v&(n_330_v&m4_v))));
  assign n_1697_v = ~((n_1618_v|(_t2_v&(n_220_v&m3_v))|(_t3_v&(n_330_v&m4_v))));
  assign n_1692_v = ~(((_t2_v&(n_271_v&m4_v))|(_t3_v&(n_220_v&m3_v))));
  assign n_1691_v = ~((_t4_v&(n_458_v&m3_v)));
  assign n_1699_v = ~(((n_1594_v|n_612_v)&(n_622_v&n_1678_v)));
  assign n_1694_v = ~(((n_271_v&m3_v)&(_t2_v|(_t4_v&n_449_v))));
  assign n_1679_v = ~(n_1668_v);
  assign n_1678_v = ~((n_1461_v&n_612_v));
  assign n_1688_v = ~(n_1486_v);
  assign n_1693_v = ~((n_542_v&n_1486_v));
  assign n_1673_v = ~(n_1682_v);
  assign n_1696_v = ~(n_1681_v);
  assign n_1710_v = ~((n_449_v&n_618_v));
  assign n_1762_v = ~((n_582_v|v(clk_v)));
  assign n_1758_v = ~((n_1704_v|v(clk_v)));
  assign n_1749_v = ~((n_609_v|n_594_v));
  assign n_1750_v = ~((n_605_v|n_594_v));
  assign n_1751_v = ~((n_605_v|n_1446_v));
  assign n_1752_v = ~((n_609_v|n_1446_v));
  assign n_1683_v = ~(n_1724_v);
  assign n_1755_v = ~((n_1678_v|v(clk_v)));
  assign n_1672_v = ~(n_1700_v);
  assign n_1759_v = ~((n_1619_v|v(clk_v)));
  assign n_1764_v = ~(n_1718_v);
  assign n_1756_v = ~(n_1721_v);
  assign n_1763_v = ~((v(clk_v)|n_1729_v));
  assign n_1757_v = ~((v(clk_v)|n_1726_v));
  assign n_1766_v = ~(n_1710_v);
  assign n_1761_v = ~((n_1734_v&m6_v));
  assign n_1723_v = ~(n_1735_v);
  assign n_1760_v = ~(m6_v);
  assign n_1765_v = ~(n_619_v);
  assign n_1790_v = ~((v(clk_v)|n_649_v));
  assign n_1769_v = ~(n_1764_v);
  assign n_1732_v = ~(n_1782_v);
  assign n_1784_v = ~(n_1831_v);
  assign n_1789_v = ~((n_1778_v&n_1761_v));
  assign n_1787_v = ~((n_644_v|v(clk_v)));
  assign n_1775_v = ~((n_1754_v&n_756_v));
  assign n_1794_v = ~((v(clk_v)|n_1780_v));
  assign n_1793_v = ~((n_638_v|v(clk_v)));
  assign n_1792_v = ~(n_686_v);
  assign n_1791_v = ~(n_1775_v);
  assign n_1786_v = ~(n_1696_v);
  assign n_1788_v = ~(n_573_v);
  assign n_1806_v = ~(v(n_1783_v));
  assign n_1801_v = ~(n_1756_v);
  assign n_1802_v = ~((n_612_v&n_1496_v));
  assign n_1805_v = ~(n_1460_v);
  assign n_1808_v = ~(n_830_v);
  assign n_1778_v = ~(v(n_696_v));
  assign n_1813_v = ~(n_1810_v);
  assign n_1839_v = ~(v(n_701_v));
  assign n_1860_v = ~((n_618_v&(n_449_v&n_1749_v)));
  assign n_1859_v = ~((n_352_v&(n_1809_v&n_819_v)));
  assign n_1811_v = ~(n_767_v);
  assign n_1838_v = ~((n_1855_v|n_692_v));
  assign n_1833_v = ~(n_704_v);
  assign n_1862_v = ~(n_1778_v);
  assign n_1858_v = ~(n_711_v);
  assign n_1857_v = ~(n_449_v);
  assign n_1812_v = ~((n_1802_v|v(clk_v)));
  assign n_1855_v = ~((v(n_708_v)|n_692_v));
  assign n_1882_v = ~((v(n_715_v)|n_692_v));
  assign n_1911_v = ~((n_352_v&(n_1864_v&n_762_v)));
  assign n_1904_v = ~(n_827_v);
  assign n_1885_v = ~(n_719_v);
  assign n_1905_v = ~((n_692_v|n_1882_v));
  assign n_1964_v = ~((n_1861_v|v(clk_v)));
  assign n_1908_v = ~(n_682_v);
  assign n_1933_v = ~((v(n_687_v)|n_648_v));
  assign n_1930_v = ~((n_720_v|v(clk_v)));
  assign n_1944_v = ~(v(n_816_v));
  assign n_1959_v = ~(n_768_v);
  assign n_1943_v = ~(n_764_v);
  assign n_1932_v = ~(n_1860_v);
  assign n_1961_v = ~(n_724_v);
  assign n_1962_v = ~(n_1789_v);
  assign n_1940_v = ~((n_1960_v|n_692_v));
  assign n_1935_v = ~(n_741_v);
  assign n_1913_v = ~((n_165_v|n_733_v));
  assign n_1965_v = ~((n_165_v|n_751_v));
  assign n_1960_v = ~((v(n_745_v)|n_692_v));
  assign n_1987_v = ~((v(n_753_v)|n_692_v));
  assign n_1989_v = ~(n_642_v);
  assign n_1991_v = ~(n_761_v);
  assign n_2010_v = ~((n_692_v|n_1987_v));
  assign n_2011_v = ~(n_682_v);
  assign n_2017_v = ~(n_610_v);
  assign n_2015_v = ~(v(db6_v));
  assign n_2016_v = ~((n_133_v|n_82_v));
  assign n_2043_v = ~(n_757_v);
  assign n_2061_v = ~(n_515_v);
  assign n_2041_v = ~((n_2059_v|n_692_v));
  assign n_2036_v = ~(n_780_v);
  assign n_2063_v = ~(n_768_v);
  assign n_2064_v = ~(n_1859_v);
  assign n_2062_v = ~(n_765_v);
  assign n_2112_v = ~((n_1572_v|v(clk_v)));
  assign n_2111_v = ~((n_1791_v|v(clk_v)));
  assign n_2066_v = ~(n_764_v);
  assign n_2109_v = ~((n_756_v|v(clk_v)));
  assign n_2059_v = ~((v(n_785_v)|n_692_v));
  assign n_2090_v = ~(n_734_v);
  assign n_2110_v = ~(n_747_v);
  assign n_2083_v = ~((v(n_799_v)|n_692_v));
  assign n_2084_v = ~(n_1911_v);
  assign n_2115_v = ~(n_747_v);
  assign n_2087_v = ~(n_801_v);
  assign n_2108_v = ~((n_692_v|n_2083_v));
  assign n_2140_v = ~((n_2156_v|n_692_v));
  assign n_2136_v = ~(n_812_v);
  assign n_2156_v = ~((v(n_834_v)|n_692_v));
  assign n_2188_v = ~(n_2161_v);
  assign n_2162_v = ~((v(n_847_v)|n_692_v));
  assign n_2181_v = ~((v(n_837_v)|n_603_v));
  assign n_2193_v = ~(n_2217_v);
  assign n_2192_v = ~(n_2189_v);
  assign n_2210_v = ~((v(n_486_v)&(v(n_485_v)&v(n_480_v))));
  assign n_2213_v = ~(n_829_v);
  assign n_2219_v = ~(((v(n_754_v)&(n_844_v&n_2186_v))|((n_844_v|n_2186_v|v(n_754_v))&(n_855_v|n_828_v))));
  assign n_2185_v = ~(n_853_v);
  assign n_2215_v = ~((n_692_v|n_2162_v));
  assign n_2212_v = ~(n_865_v);
  assign n_2189_v = ~(v(n_850_v));
  assign n_2216_v = ~((n_2181_v|n_603_v));
  assign n_2214_v = ~((n_859_v|n_165_v));
  assign n_2217_v = ~(v(n_845_v));
  assign n_2223_v = ~(((n_747_v&((n_2193_v&n_757_v)|(n_2217_v&n_823_v)))|(n_824_v&((n_2224_v&n_823_v)|(n_2255_v&n_757_v)))));
  assign n_2218_v = ~(v(n_2211_v));
  assign n_2224_v = ~(v(n_867_v));
  assign n_2226_v = ~(n_868_v);
  assign n_2191_v = ~(n_2212_v);
  assign n_2227_v = ~((n_883_v&(v(n_480_v)&v(n_485_v))));
  assign n_2228_v = ~((n_603_v|n_2231_v));
  assign n_2230_v = ~(n_2223_v);
  assign n_2247_v = ~(n_2219_v);
  assign n_2231_v = ~((n_603_v|v(n_852_v)));
  assign n_2256_v = ~(n_2226_v);
  assign n_2254_v = ~((n_2274_v|n_693_v));
  assign n_2250_v = ~(n_873_v);
  assign n_2255_v = ~(n_2224_v);
  assign n_2229_v = ~((n_872_v|n_165_v));
  assign n_2273_v = ~(n_869_v);
  assign n_2272_v = ~(n_2276_v);
  assign n_2274_v = ~((v(n_880_v)|n_693_v));
  assign n_2277_v = ~(v(db5_v));
  assign n_2297_v = ~((v(n_886_v)|n_693_v));
  assign n_2300_v = ~(n_890_v);
  assign n_2321_v = ~((n_693_v|n_2297_v));
  assign n_2331_v = ~(n_2322_v);
  assign n_2326_v = ~((v(n_889_v)|n_603_v));
  assign n_2337_v = ~(n_2342_v);
  assign n_2335_v = ~(n_2332_v);
  assign n_2360_v = ~(((n_878_v&(n_896_v&n_2330_v))|((n_896_v|n_2330_v|n_878_v)&(n_904_v|n_828_v))));
  assign n_2340_v = ~(n_876_v);
  assign n_2324_v = ~(n_872_v);
  assign n_2323_v = ~((n_883_v|v(n_480_v)|n_2370_v));
  assign n_2339_v = ~(n_912_v);
  assign n_2333_v = ~(n_2323_v);
  assign n_2332_v = ~(v(n_899_v));
  assign n_2367_v = ~((n_2385_v|n_693_v));
  assign n_2363_v = ~(n_909_v);
  assign n_2341_v = ~((n_2326_v|n_603_v));
  assign n_2342_v = ~(v(n_897_v));
  assign n_2369_v = ~(((n_747_v&((n_2337_v&n_757_v)|(n_2342_v&n_823_v)))|(n_824_v&((n_2388_v&n_823_v)|(n_2399_v&n_757_v)))));
  assign n_2358_v = ~(v(n_2338_v));
  assign n_2336_v = ~(n_2324_v);
  assign n_2370_v = ~(v(n_485_v));
  assign n_2388_v = ~(v(n_918_v));
  assign n_2390_v = ~(n_920_v);
  assign n_2385_v = ~((v(n_914_v)|n_693_v));
  assign n_2334_v = ~(n_2339_v);
  assign n_2392_v = ~((n_603_v|n_2395_v));
  assign n_2391_v = ~((n_2370_v|v(n_486_v)|v(n_480_v)));
  assign n_2393_v = ~(n_2369_v);
  assign n_2389_v = ~((n_82_v|n_133_v));
  assign n_2397_v = ~(n_2360_v);
  assign n_2395_v = ~((n_603_v|v(n_903_v)));
  assign n_2400_v = ~(n_2390_v);
  assign n_2398_v = ~(n_2391_v);
  assign n_2399_v = ~(n_2388_v);
  assign n_2417_v = ~((v(n_923_v)|n_693_v));
  assign n_2426_v = ~(n_919_v);
  assign n_2423_v = ~(n_2443_v);
  assign n_2425_v = ~((n_133_v|n_82_v));
  assign n_2420_v = ~(n_927_v);
  assign n_2444_v = ~((n_693_v|n_2417_v));
  assign n_2445_v = ~(n_2447_v);
  assign n_2447_v = ~(n_930_v);
  assign n_2471_v = ~((n_2490_v|n_693_v));
  assign n_2467_v = ~(n_938_v);
  assign n_2497_v = ~(n_2474_v);
  assign n_2491_v = ~((v(n_937_v)|n_603_v));
  assign n_2501_v = ~(n_2498_v);
  assign n_2502_v = ~(n_2509_v);
  assign n_2490_v = ~((v(n_949_v)|n_693_v));
  assign n_2503_v = ~(v(n_908_v));
  assign n_2511_v = ~(((n_925_v&(n_943_v&n_2496_v))|((n_943_v|n_2496_v|n_925_v)&(n_952_v|n_828_v))));
  assign n_2475_v = ~((v(n_485_v)|n_883_v|n_2530_v));
  assign n_2499_v = ~(n_2475_v);
  assign n_2505_v = ~(n_960_v);
  assign n_2498_v = ~(v(n_947_v));
  assign n_2528_v = ~((v(n_959_v)|n_693_v));
  assign n_2508_v = ~((n_2491_v|n_603_v));
  assign n_2509_v = ~(v(n_944_v));
  assign n_2531_v = ~(((n_747_v&((n_2502_v&n_757_v)|(n_2509_v&n_823_v)))|(n_824_v&((n_2554_v&n_823_v)|(n_2567_v&n_757_v)))));
  assign n_2510_v = ~(v(n_2504_v));
  assign n_2535_v = ~(v(db3_v));
  assign n_2530_v = ~(v(n_480_v));
  assign n_2533_v = ~(n_962_v);
  assign n_2555_v = ~((n_693_v|n_2528_v));
  assign n_2556_v = ~(n_968_v);
  assign n_2554_v = ~(v(n_966_v));
  assign n_2500_v = ~(n_2505_v);
  assign n_2558_v = ~((n_603_v|n_2561_v));
  assign n_2557_v = ~((n_2530_v|v(n_486_v)|v(n_485_v)));
  assign n_2560_v = ~(n_2531_v);
  assign n_2563_v = ~(n_2511_v);
  assign n_2561_v = ~((n_603_v|v(n_951_v)));
  assign n_2566_v = ~(n_2556_v);
  assign n_2565_v = ~(v(n_956_v));
  assign n_2564_v = ~(n_2557_v);
  assign n_2567_v = ~(n_2554_v);
  assign n_2568_v = ~((n_165_v|n_930_v));
  assign n_2571_v = ~(n_967_v);
  assign n_2570_v = ~(n_2595_v);
  assign n_2594_v = ~((n_2611_v|n_693_v));
  assign n_2590_v = ~(n_975_v);
  assign n_2611_v = ~((v(n_980_v)|n_693_v));
  assign n_2613_v = ~((n_165_v|n_978_v));
  assign n_2634_v = ~((v(n_985_v)|n_693_v));
  assign n_2661_v = ~(n_2635_v);
  assign n_2641_v = ~((v(n_983_v)|n_603_v));
  assign n_2666_v = ~(n_2673_v);
  assign n_2667_v = ~(n_2662_v);
  assign n_2637_v = ~(n_990_v);
  assign n_2665_v = ~((n_693_v|n_2634_v));
  assign n_2638_v = ~((v(n_485_v)|n_883_v|v(n_480_v)));
  assign n_2670_v = ~(n_2658_v);
  assign n_2669_v = ~((n_133_v|n_82_v));
  assign n_2676_v = ~(((n_767_v&(n_989_v&n_2659_v))|((n_989_v|n_2659_v|n_767_v)&(n_997_v|n_828_v))));
  assign n_2663_v = ~(n_2638_v);
  assign n_2668_v = ~(n_1002_v);
  assign n_2662_v = ~(v(n_993_v));
  assign n_2672_v = ~((n_2641_v|n_603_v));
  assign n_2677_v = ~(n_2679_v);
  assign n_2673_v = ~(v(n_988_v));
  assign n_2678_v = ~(((n_747_v&((n_2666_v&n_757_v)|(n_2673_v&n_823_v)))|(n_824_v&((n_2680_v&n_823_v)|(n_2690_v&n_757_v)))));
  assign n_2675_v = ~(v(n_816_v));
  assign n_2679_v = ~(n_1000_v);
  assign n_2681_v = ~((v(n_480_v)|v(n_485_v)|v(n_486_v)));
  assign n_2680_v = ~(v(n_1005_v));
  assign n_2682_v = ~(n_1007_v);
  assign n_2664_v = ~(n_2668_v);
  assign n_2684_v = ~((n_603_v|n_2685_v));
  assign n_2685_v = ~((n_603_v|v(n_995_v)));
  assign n_2683_v = ~(n_2678_v);
  assign n_2686_v = ~(n_2676_v);
  assign n_2687_v = ~(n_2681_v);
  assign n_2688_v = ~(v(n_1001_v));
  assign n_2691_v = ~(n_2682_v);
  assign n_2690_v = ~(n_2680_v);
  assign n_2693_v = ~(n_1006_v);
  assign n_2692_v = ~(n_2694_v);
  assign n_2697_v = ~((n_165_v|n_1011_v));
  assign n_2699_v = ~(v(n_486_v));
  assign n_2707_v = ~((n_165_v|n_1000_v));
  assign n_2709_v = ~((n_1013_v|n_627_v));
  assign n_2716_v = ~((n_1015_v|n_627_v));
  assign n_2717_v = ~((n_1016_v|n_627_v));
  assign n_2718_v = ~((n_1019_v|n_627_v));
  assign n_2726_v = ~((n_627_v|v(n_2705_v)));
  assign n_2714_v = ~((n_627_v|n_1025_v));
  assign n_2724_v = ~(n_1025_v);
  assign n_2737_v = ~(n_1013_v);
  assign n_2738_v = ~(n_1015_v);
  assign n_2739_v = ~(n_1016_v);
  assign n_2740_v = ~(n_1019_v);
  assign n_2749_v = ~((n_627_v|v(n_1020_v)));
  assign n_2750_v = ~((v(n_1014_v)|n_627_v));
  assign n_2752_v = ~((n_627_v|v(n_1017_v)));
  assign n_2753_v = ~((v(n_1018_v)|n_627_v));

  spice_mux_3 mux_12004(eclk, ereset, n_2037_v,n_2018_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_2617_v), n_792_v);
  spice_mux_2 mux_12005(eclk, ereset, n_1069_v,v(n_1072_v), 1'b1,1'b0, n_1042_v);
  spice_mux_2 mux_12006(eclk, ereset, n_1108_v,(v(n_81_v)|n_69_v), 1'b1,1'b0, n_1039_v);
  spice_mux_2 mux_12007(eclk, ereset, n_1039_v,n_1040_v, 1'b1,1'b0, _rd_v);
  spice_mux_2 mux_12008(eclk, ereset, n_1249_v,v(n_185_v), 1'b1,1'b0, n_95_v);
  spice_mux_2 mux_12009(eclk, ereset, n_1346_v,v(n_216_v), 1'b1,1'b0, n_371_v);
  spice_mux_3 mux_12010(eclk, ereset, n_781_v,n_782_v,n_1798_v, 1'b1,1'b0,v(n_791_v), n_3421_v);
  spice_mux_3 mux_12011(eclk, ereset, n_2036_v,n_780_v,n_678_v, 1'b1,1'b0,v(n_785_v), n_3420_v);
  spice_mux_2 mux_12012(eclk, ereset, n_1717_v,n_1695_v, 1'b1,1'b0, n_608_v);
  spice_mux_2 mux_12013(eclk, ereset, v(n_1498_v),(v(n_1466_v)&n_431_v), 1'b1,1'b0, n_220_v);
  spice_mux_3 mux_12014(eclk, ereset, n_706_v,n_705_v,n_1798_v, 1'b1,1'b0,v(n_703_v), n_3366_v);
  spice_mux_3 mux_12015(eclk, ereset, n_911_v,n_910_v,n_1798_v, 1'b1,1'b0,v(n_907_v), n_3493_v);
  spice_mux_2 mux_12016(eclk, ereset, n_2043_v,n_757_v, 1'b1,1'b0, n_823_v);
  spice_mux_3 mux_12017(eclk, ereset, n_823_v,n_757_v,n_551_v, 1'b1,1'b0,v(n_528_v), n_794_v);
  spice_mux_3 mux_12018(eclk, ereset, n_909_v,n_2363_v,n_652_v, 1'b1,1'b0,v(n_906_v), n_3494_v);
  spice_mux_3 mux_12019(eclk, ereset, n_704_v,n_1833_v,n_678_v, 1'b1,1'b0,v(n_702_v), n_3367_v);
  spice_mux_2 mux_12020(eclk, ereset, n_1203_v,(n_123_v|n_165_v), 1'b1,1'b0, n_170_v);
  spice_mux_2 mux_12021(eclk, ereset, n_1241_v,v(n_1225_v), 1'b1,1'b0, m4_v);
  spice_mux_2 mux_12022(eclk, ereset, n_1359_v,n_373_v, 1'b1,1'b0, n_1358_v);
  spice_mux_2 mux_12023(eclk, ereset, n_1104_v,(v(n_86_v)|n_69_v), 1'b1,1'b0, n_100_v);
  spice_mux_2 mux_12024(eclk, ereset, n_100_v,n_1042_v, 1'b1,1'b0, _mreq_v);
  spice_mux_2 mux_12025(eclk, ereset, n_1372_v,(n_358_v|n_165_v), 1'b1,1'b0, n_383_v);
  spice_mux_3 mux_12026(eclk, ereset, n_1362_v,n_1363_v,n_87_v, 1'b1,1'b0,v(n_370_v), n_2937_v);
  spice_mux_2 mux_12027(eclk, ereset, n_373_v,n_1359_v, 1'b1,1'b0, n_375_v);
  spice_mux_2 mux_12028(eclk, ereset, n_1156_v,n_1155_v, 1'b1,1'b0, n_99_v);
  spice_mux_2 mux_12029(eclk, ereset, n_1330_v,(n_195_v|n_165_v), 1'b1,1'b0, n_250_v);
  spice_mux_2 mux_12030(eclk, ereset, n_1309_v,n_226_v, 1'b1,1'b0, n_254_v);
  spice_mux_2 mux_12031(eclk, ereset, n_1505_v,n_1504_v, 1'b1,1'b0, n_588_v);
  spice_mux_3 mux_12032(eclk, ereset, n_1834_v,n_1776_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_689_v), n_3372_v);
  spice_mux_2 mux_12033(eclk, ereset, n_1510_v,(n_487_v|n_87_v), 1'b1,1'b0, n_1507_v);
  spice_mux_3 mux_12034(eclk, ereset, n_2364_v,n_2343_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_2704_v), n_2396_v);
  spice_mux_2 mux_12035(eclk, ereset, n_1801_v,n_1756_v, 1'b1,1'b0, n_795_v);
  spice_mux_3 mux_12036(eclk, ereset, n_705_v,n_706_v,n_1798_v, 1'b1,1'b0,v(n_713_v), n_3375_v);
  spice_mux_3 mux_12037(eclk, ereset, n_800_v,n_805_v,n_1798_v, 1'b1,1'b0,v(n_798_v), n_3424_v);
  spice_mux_3 mux_12038(eclk, ereset, n_910_v,n_911_v,n_1798_v, 1'b1,1'b0,v(n_917_v), n_3499_v);
  spice_mux_3 mux_12039(eclk, ereset, n_2363_v,n_909_v,n_652_v, 1'b1,1'b0,v(n_914_v), n_3498_v);
  spice_mux_3 mux_12040(eclk, ereset, n_1833_v,n_704_v,n_678_v, 1'b1,1'b0,v(n_708_v), n_3374_v);
  spice_mux_2 mux_12041(eclk, ereset, n_1247_v,v(n_1221_v), 1'b1,1'b0, m5_v);
  spice_mux_2 mux_12042(eclk, ereset, n_1312_v,n_1254_v, 1'b1,1'b0, n_192_v);
  spice_mux_2 mux_12043(eclk, ereset, n_1644_v,n_1630_v, 1'b1,1'b0, n_600_v);
  spice_mux_2 mux_12044(eclk, ereset, n_1651_v,n_1650_v, 1'b1,1'b0, n_602_v);
  spice_mux_2 mux_12045(eclk, ereset, n_1365_v,n_376_v, 1'b1,1'b0, n_1364_v);
  spice_mux_2 mux_12046(eclk, ereset, n_1511_v,n_493_v, 1'b1,1'b0, n_465_v);
  spice_mux_3 mux_12047(eclk, ereset, n_2084_v,n_1911_v,n_795_v, 1'b1,1'b0,v(n_528_v), n_3415_v);
  spice_mux_2 mux_12048(eclk, ereset, n_1318_v,n_252_v, 1'b1,1'b0, n_177_v);
  spice_mux_3 mux_12049(eclk, ereset, n_829_v,n_686_v,n_551_v, 1'b1,1'b0,v(n_526_v), n_3412_v);
  spice_mux_3 mux_12050(eclk, ereset, n_2061_v,n_515_v,n_551_v, 1'b1,1'b0,v(n_716_v), n_3416_v);
  spice_mux_3 mux_12051(eclk, ereset, n_2084_v,n_1911_v,n_795_v, 1'b1,1'b0,v(n_526_v), n_3411_v);
  spice_mux_3 mux_12052(eclk, ereset, n_2087_v,n_801_v,n_678_v, 1'b1,1'b0,v(n_799_v), n_3426_v);
  spice_mux_3 mux_12053(eclk, ereset, n_2063_v,n_768_v,n_551_v, 1'b1,1'b0,v(n_525_v), n_3407_v);
  spice_mux_3 mux_12054(eclk, ereset, n_2086_v,n_2088_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_1009_v), n_797_v);
  spice_mux_3 mux_12055(eclk, ereset, n_2066_v,n_764_v,n_551_v, 1'b1,1'b0,v(n_545_v), n_3414_v);
  spice_mux_2 mux_12056(eclk, ereset, n_2386_v,(v(n_2320_v)|n_627_v), 1'b1,1'b0, n_2421_v);
  spice_mux_2 mux_12057(eclk, ereset, n_2117_v,(n_627_v|v(n_2116_v)), 1'b1,1'b0, n_2091_v);
  spice_mux_2 mux_12058(eclk, ereset, n_2091_v,n_2044_v, 1'b1,1'b0, ab2_v);
  spice_mux_2 mux_12059(eclk, ereset, n_1514_v,n_1513_v, 1'b1,1'b0, n_589_v);
  spice_mux_2 mux_12060(eclk, ereset, n_924_v,(n_825_v|n_904_v), 1'b1,1'b0, n_925_v);
  spice_mux_3 mux_12061(eclk, ereset, n_2388_v,n_2399_v,n_574_v, 1'b1,1'b0,v(n_903_v), n_3509_v);
  spice_mux_2 mux_12062(eclk, ereset, n_376_v,n_1365_v, 1'b1,1'b0, n_378_v);
  spice_mux_3 mux_12063(eclk, ereset, n_2064_v,n_1859_v,n_795_v, 1'b1,1'b0,v(n_716_v), n_3413_v);
  spice_mux_3 mux_12064(eclk, ereset, n_2064_v,n_1859_v,n_795_v, 1'b1,1'b0,v(n_790_v), n_3409_v);
  spice_mux_2 mux_12065(eclk, ereset, n_1658_v,n_578_v, 1'b1,1'b0, n_1674_v);
  spice_mux_3 mux_12066(eclk, ereset, n_2390_v,n_2400_v,n_552_v, 1'b1,1'b0,v(n_903_v), n_3511_v);
  spice_mux_3 mux_12067(eclk, ereset, n_926_v,n_931_v,n_1798_v, 1'b1,1'b0,v(n_922_v), n_3506_v);
  spice_mux_3 mux_12068(eclk, ereset, n_2062_v,n_765_v,n_551_v, 1'b1,1'b0,v(n_779_v), n_3408_v);
  spice_mux_2 mux_12069(eclk, ereset, n_1317_v,n_1299_v, 1'b1,1'b0, n_267_v);
  spice_mux_2 mux_12070(eclk, ereset, n_1661_v,n_598_v, 1'b1,1'b0, n_750_v);
  spice_mux_3 mux_12071(eclk, ereset, n_788_v,n_786_v,n_87_v, 1'b1,1'b0,v(n_380_v), n_3428_v);
  spice_mux_3 mux_12072(eclk, ereset, n_1408_v,n_1409_v,n_87_v, 1'b1,1'b0,v(n_412_v), n_2971_v);
  spice_mux_2 mux_12073(eclk, ereset, n_1665_v,(v(n_562_v)|(n_1609_v&v(clk_v))), 1'b1,1'b0, n_627_v);
  spice_mux_2 mux_12074(eclk, ereset, n_2109_v,(n_756_v|v(clk_v)), 1'b1,1'b0, n_822_v);
  spice_mux_2 mux_12075(eclk, ereset, n_2111_v,(n_1791_v|v(clk_v)), 1'b1,1'b0, n_821_v);
  spice_mux_2 mux_12076(eclk, ereset, n_1316_v,n_1297_v, 1'b1,1'b0, n_263_v);
  spice_mux_2 mux_12077(eclk, ereset, n_1369_v,n_379_v, 1'b1,1'b0, n_1368_v);
  spice_mux_2 mux_12078(eclk, ereset, n_2112_v,(n_1572_v|v(clk_v)), 1'b1,1'b0, n_820_v);
  spice_mux_2 mux_12079(eclk, ereset, n_1202_v,(v(clk_v)|n_1195_v), 1'b1,1'b0, n_133_v);
  spice_mux_3 mux_12080(eclk, ereset, n_2420_v,n_927_v,n_652_v, 1'b1,1'b0,v(n_923_v), n_3508_v);
  spice_mux_3 mux_12081(eclk, ereset, n_2419_v,n_2422_v,(v(clk_v)&n_393_v), 1'b1,1'b0,v(n_2705_v), n_921_v);
  spice_mux_2 mux_12082(eclk, ereset, n_2393_v,n_2369_v, 1'b1,1'b0, n_2330_v);
  spice_mux_3 mux_12083(eclk, ereset, n_2398_v,n_2391_v,n_553_v, 1'b1,1'b0,v(n_903_v), n_3513_v);
  spice_mux_2 mux_12084(eclk, ereset, n_379_v,n_1369_v, 1'b1,1'b0, n_1371_v);
  spice_mux_3 mux_12085(eclk, ereset, n_805_v,n_800_v,n_1798_v, 1'b1,1'b0,v(n_806_v), n_3429_v);
  spice_mux_2 mux_12086(eclk, ereset, n_1679_v,n_1668_v, 1'b1,1'b0, n_603_v);
  spice_mux_3 mux_12087(eclk, ereset, n_801_v,n_2087_v,n_678_v, 1'b1,1'b0,v(n_807_v), n_3430_v);
  spice_mux_2 mux_12088(eclk, ereset, n_2110_v,n_747_v, 1'b1,1'b0, n_831_v);
  spice_mux_2 mux_12089(eclk, ereset, n_1418_v,v(n_408_v), 1'b1,1'b0, n_436_v);
  spice_mux_2 mux_12090(eclk, ereset, n_1762_v,(n_582_v|v(clk_v)), 1'b1,1'b0, n_832_v);
  spice_mux_3 mux_12091(eclk, ereset, n_832_v,v(clk_v),n_604_v, 1'b1,n_2400_v,v(n_903_v), n_920_v);
  spice_mux_2 mux_12092(eclk, ereset, n_2426_v,n_919_v, 1'b1,1'b0, n_896_v);
  spice_mux_2 mux_12093(eclk, ereset, n_2115_v,n_747_v, 1'b1,1'b0, n_824_v);
  spice_mux_2 mux_12094(eclk, ereset, n_1680_v,(n_1654_v|v(clk_v)), 1'b1,1'b0, n_604_v);
  spice_mux_3 mux_12095(eclk, ereset, n_718_v,n_725_v,n_1798_v, 1'b1,1'b0,v(n_714_v), n_3381_v);
  spice_mux_2 mux_12096(eclk, ereset, n_1965_v,(n_751_v|n_165_v), 1'b1,1'b0, n_733_v);
  spice_mux_3 mux_12097(eclk, ereset, n_931_v,n_926_v,n_1798_v, 1'b1,1'b0,v(n_933_v), n_3514_v);
  spice_mux_3 mux_12098(eclk, ereset, n_927_v,n_2420_v,n_652_v, 1'b1,1'b0,v(n_934_v), n_3515_v);
  spice_mux_2 mux_12099(eclk, ereset, n_2421_v,n_2492_v, 1'b1,1'b0, ab3_v);
  spice_mux_2 mux_12100(eclk, ereset, n_1374_v,n_382_v, 1'b1,1'b0, n_1373_v);
  spice_mux_2 mux_12101(eclk, ereset, n_1270_v,n_1272_v, 1'b1,1'b0, n_103_v);
  spice_mux_2 mux_12102(eclk, ereset, n_371_v,n_1385_v, 1'b1,1'b0, _m1_v);
  spice_mux_2 mux_12103(eclk, ereset, n_386_v,(n_389_v|n_65_v), 1'b1,1'b0, n_107_v);
  spice_mux_2 mux_12104(eclk, ereset, n_382_v,n_1374_v, 1'b1,1'b0, n_1377_v);
  spice_mux_2 mux_12105(eclk, ereset, n_1056_v,(n_1048_v|n_60_v), 1'b1,1'b0, n_59_v);
  spice_mux_2 mux_12106(eclk, ereset, n_1328_v,n_1334_v, 1'b1,1'b0, n_126_v);
  spice_mux_3 mux_12107(eclk, ereset, n_1885_v,n_719_v,n_678_v, 1'b1,1'b0,v(n_715_v), n_3385_v);
  spice_mux_3 mux_12108(eclk, ereset, n_1883_v,n_1886_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_723_v), n_3383_v);
  spice_mux_2 mux_12109(eclk, ereset, n_1154_v,(v(n_92_v)|n_105_v), 1'b1,1'b0, _t1_v);
  spice_mux_2 mux_12110(eclk, ereset, n_1063_v,n_108_v, 1'b1,1'b0, n_1035_v);
  spice_mux_2 mux_12111(eclk, ereset, n_1035_v,n_108_v, 1'b1,1'b0, _halt_v);
  spice_mux_2 mux_12112(eclk, ereset, v(n_1332_v),v(n_241_v), 1'b1,1'b0, m6_v);
  spice_mux_2 mux_12113(eclk, ereset, n_1378_v,(n_383_v|n_165_v), 1'b1,1'b0, n_1376_v);
  spice_mux_2 mux_12114(eclk, ereset, n_1045_v,n_63_v, 1'b1,1'b0, n_64_v);
  spice_mux_2 mux_12115(eclk, ereset, n_388_v,n_1379_v, 1'b1,1'b0, n_385_v);
  spice_mux_2 mux_12116(eclk, ereset, v(n_73_v),v(n_70_v), 1'b1,1'b0, n_106_v);
  spice_mux_3 mux_12117(eclk, ereset, n_815_v,n_814_v,n_1798_v, 1'b1,1'b0,v(n_810_v), n_3432_v);
  spice_mux_3 mux_12118(eclk, ereset, n_941_v,n_939_v,n_1798_v, 1'b1,1'b0,v(n_936_v), n_3518_v);
  spice_mux_3 mux_12119(eclk, ereset, n_812_v,n_2136_v,n_678_v, 1'b1,1'b0,v(n_809_v), n_3433_v);
  spice_mux_3 mux_12120(eclk, ereset, n_938_v,n_2467_v,n_652_v, 1'b1,1'b0,v(n_935_v), n_3519_v);
  spice_mux_3 mux_12121(eclk, ereset, n_1533_v,n_514_v,n_1757_v, 1'b1,1'b0,v(n_647_v), n_502_v);
  spice_mux_3 mux_12122(eclk, ereset, n_1181_v,n_117_v,n_87_v, 1'b1,1'b0,v(n_138_v), n_2820_v);
  spice_mux_2 mux_12123(eclk, ereset, n_1381_v,(n_65_v|n_390_v), 1'b1,1'b0, n_393_v);
  spice_mux_2 mux_12124(eclk, ereset, n_1047_v,n_53_v, 1'b1,1'b0, n_54_v);
  spice_mux_3 mux_12125(eclk, ereset, n_1387_v,n_392_v,n_180_v, 1'b1,1'b0,n_179_v, n_247_v);
  spice_mux_3 mux_12126(eclk, ereset, n_725_v,n_718_v,n_1798_v, 1'b1,1'b0,v(n_731_v), n_3389_v);
  spice_mux_3 mux_12127(eclk, ereset, n_2445_v,n_2447_v,n_87_v, 1'b1,1'b0,v(n_480_v), n_3522_v);
  spice_mux_2 mux_12128(eclk, ereset, n_1074_v,(n_69_v|v(n_85_v)), 1'b1,1'b0, n_1038_v);
  spice_mux_3 mux_12129(eclk, ereset, n_2468_v,n_2449_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_1020_v), n_954_v);
  spice_mux_3 mux_12130(eclk, ereset, n_719_v,n_1885_v,n_678_v, 1'b1,1'b0,v(n_732_v), n_3390_v);
  spice_mux_2 mux_12131(eclk, ereset, n_1884_v,(v(n_723_v)|n_627_v), 1'b1,1'b0, n_1912_v);
  spice_mux_3 mux_12132(eclk, ereset, n_2137_v,n_2118_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_2700_v), n_2160_v);
  spice_mux_3 mux_12133(eclk, ereset, n_2499_v,n_2475_v,n_553_v, 1'b1,1'b0,v(n_937_v), n_3521_v);
  spice_mux_3 mux_12134(eclk, ereset, n_2498_v,n_2501_v,n_552_v, 1'b1,1'b0,v(n_937_v), n_3523_v);
  spice_mux_3 mux_12135(eclk, ereset, n_939_v,n_941_v,n_1798_v, 1'b1,1'b0,v(n_953_v), n_3529_v);
  spice_mux_3 mux_12136(eclk, ereset, n_2500_v,n_2505_v,n_646_v, 1'b1,1'b0,v(n_937_v), n_2494_v);
  spice_mux_3 mux_12137(eclk, ereset, n_2467_v,n_938_v,n_652_v, 1'b1,1'b0,v(n_949_v), n_3527_v);
  spice_mux_2 mux_12138(eclk, ereset, n_392_v,n_1387_v, 1'b1,1'b0, n_1386_v);
  spice_mux_2 mux_12139(eclk, ereset, n_2506_v,(n_627_v|n_905_v), 1'b1,1'b0, n_2492_v);
  spice_mux_2 mux_12140(eclk, ereset, n_1428_v,(n_165_v|n_414_v), 1'b1,1'b0, n_452_v);
  spice_mux_3 mux_12141(eclk, ereset, n_814_v,n_815_v,n_1798_v, 1'b1,1'b0,v(n_841_v), n_3436_v);
  spice_mux_3 mux_12142(eclk, ereset, n_2509_v,n_2502_v,n_574_v, 1'b1,1'b0,v(n_937_v), n_3525_v);
  spice_mux_3 mux_12143(eclk, ereset, n_2136_v,n_812_v,n_678_v, 1'b1,1'b0,v(n_834_v), n_3435_v);
  spice_mux_2 mux_12144(eclk, ereset, n_1912_v,n_1966_v, 1'b1,1'b0, ab1_v);
  spice_mux_2 mux_12145(eclk, ereset, n_1075_v,v(n_1077_v), 1'b1,1'b0, n_87_v);
  spice_mux_2 mux_12146(eclk, ereset, n_1394_v,n_397_v, 1'b1,1'b0, n_1390_v);
  spice_mux_2 mux_12147(eclk, ereset, n_1086_v,n_1067_v, 1'b1,1'b0, n_83_v);
  spice_mux_2 mux_12148(eclk, ereset, n_1430_v,n_327_v, 1'b1,1'b0, n_1440_v);
  spice_mux_2 mux_12149(eclk, ereset, n_1440_v,n_1462_v, 1'b1,1'b0, _rfsh_v);
  spice_mux_2 mux_12150(eclk, ereset, n_1186_v,n_184_v, 1'b1,1'b0, n_101_v);
  spice_mux_2 mux_12151(eclk, ereset, n_1088_v,n_64_v, 1'b1,1'b0, n_1036_v);
  spice_mux_2 mux_12152(eclk, ereset, n_1071_v,v(n_77_v), 1'b1,1'b0, n_90_v);
  spice_mux_2 mux_12153(eclk, ereset, n_1434_v,n_387_v, 1'b1,1'b0, n_456_v);
  spice_mux_2 mux_12154(eclk, ereset, n_1913_v,(n_733_v|n_165_v), 1'b1,1'b0, n_1753_v);
  spice_mux_3 mux_12155(eclk, ereset, n_961_v,n_965_v,n_1798_v, 1'b1,1'b0,v(n_958_v), n_3534_v);
  spice_mux_2 mux_12156(eclk, ereset, n_1117_v,(v(n_120_v)|n_69_v), 1'b1,1'b0, n_1058_v);
  spice_mux_2 mux_12157(eclk, ereset, n_1280_v,n_182_v, 1'b1,1'b0, n_228_v);
  spice_mux_2 mux_12158(eclk, ereset, n_1216_v,(v(n_118_v)|v(n_176_v)), 1'b1,1'b0, _t3_v);
  spice_mux_3 mux_12159(eclk, ereset, n_851_v,n_858_v,n_1798_v, 1'b1,1'b0,v(n_846_v), n_3441_v);
  spice_mux_2 mux_12160(eclk, ereset, n_1441_v,(n_452_v|n_165_v), 1'b1,1'b0, n_1439_v);
  spice_mux_3 mux_12161(eclk, ereset, n_1288_v,n_1290_v,n_87_v, 1'b1,1'b0,v(n_196_v), n_2882_v);
  spice_mux_2 mux_12162(eclk, ereset, n_1058_v,n_119_v, 1'b1,1'b0, _wr_v);
  spice_mux_2 mux_12163(eclk, ereset, n_1118_v,v(n_1126_v), 1'b1,1'b0, n_108_v);
  spice_mux_2 mux_12164(eclk, ereset, n_1455_v,n_424_v, 1'b1,1'b0, n_395_v);
  spice_mux_3 mux_12165(eclk, ereset, n_2533_v,n_962_v,n_652_v, 1'b1,1'b0,v(n_959_v), n_3536_v);
  spice_mux_2 mux_12166(eclk, ereset, n_1286_v,(n_1251_v|v(clk_v)), 1'b1,1'b0, n_204_v);
  spice_mux_3 mux_12167(eclk, ereset, n_743_v,n_742_v,n_1798_v, 1'b1,1'b0,v(n_739_v), n_3392_v);
  spice_mux_3 mux_12168(eclk, ereset, n_2532_v,n_2534_v,(v(clk_v)&n_393_v), 1'b1,1'b0,v(n_1014_v), n_957_v);
  spice_mux_3 mux_12169(eclk, ereset, n_2185_v,n_853_v,n_678_v, 1'b1,1'b0,v(n_847_v), n_3443_v);
  spice_mux_3 mux_12170(eclk, ereset, n_2182_v,n_2187_v,(v(clk_v)&n_393_v), 1'b1,1'b0,v(n_2701_v), n_2163_v);
  spice_mux_3 mux_12171(eclk, ereset, n_2189_v,n_2192_v,n_552_v, 1'b1,1'b0,v(n_837_v), n_3440_v);
  spice_mux_3 mux_12172(eclk, ereset, n_741_v,n_1935_v,n_678_v, 1'b1,1'b0,v(n_738_v), n_3393_v);
  spice_mux_3 mux_12173(eclk, ereset, n_2191_v,n_2212_v,n_646_v, 1'b1,1'b0,v(n_837_v), n_2184_v);
  spice_mux_2 mux_12174(eclk, ereset, n_1932_v,n_1860_v, 1'b1,1'b0, n_734_v);
  spice_mux_2 mux_12175(eclk, ereset, n_1113_v,v(n_128_v), 1'b1,1'b0, n_119_v);
  spice_mux_3 mux_12176(eclk, ereset, n_2210_v,n_838_v,n_553_v, 1'b1,1'b0,v(n_837_v), n_3439_v);
  spice_mux_2 mux_12177(eclk, ereset, n_1120_v,(n_121_v|v(clk_v)), 1'b1,1'b0, n_122_v);
  spice_mux_2 mux_12178(eclk, ereset, n_1804_v,(n_627_v|v(n_689_v)), 1'b1,1'b0, n_1748_v);
  spice_mux_2 mux_12179(eclk, ereset, n_1748_v,(n_641_v|v(n_1709_v)), 1'b1,1'b0, ab0_v);
  spice_mux_3 mux_12180(eclk, ereset, n_2217_v,n_2193_v,n_574_v, 1'b1,1'b0,v(n_837_v), n_3444_v);
  spice_mux_2 mux_12181(eclk, ereset, n_2214_v,(n_165_v|n_859_v), 1'b1,1'b0, n_2158_v);
  spice_mux_2 mux_12182(eclk, ereset, n_1295_v,v(n_1271_v), 1'b1,1'b0, _t4_v);
  spice_mux_3 mux_12183(eclk, ereset, n_965_v,n_961_v,n_1798_v, 1'b1,1'b0,v(n_969_v), n_3541_v);
  spice_mux_2 mux_12184(eclk, ereset, n_64_v,n_1036_v, 1'b1,1'b0, _busak_v);
  spice_mux_2 mux_12185(eclk, ereset, n_1214_v,(n_178_v|n_204_v), 1'b1,1'b0, n_142_v);
  spice_mux_2 mux_12186(eclk, ereset, n_2553_v,(n_971_v|n_627_v), 1'b1,1'b0, n_2569_v);
  spice_mux_3 mux_12187(eclk, ereset, n_962_v,n_2533_v,n_652_v, 1'b1,1'b0,v(n_970_v), n_3542_v);
  spice_mux_2 mux_12188(eclk, ereset, n_972_v,(n_825_v|n_952_v), 1'b1,1'b0, n_767_v);
  spice_mux_2 mux_12189(eclk, ereset, n_1065_v,n_1057_v, 1'b1,1'b0, n_69_v);
  spice_mux_2 mux_12190(eclk, ereset, n_1933_v,(n_648_v|v(n_687_v)), 1'b1,1'b0, n_747_v);
  spice_mux_3 mux_12191(eclk, ereset, n_2554_v,n_2567_v,n_574_v, 1'b1,1'b0,v(n_951_v), n_3546_v);
  spice_mux_2 mux_12192(eclk, ereset, n_1193_v,v(n_149_v), 1'b1,1'b0, n_188_v);
  spice_mux_2 mux_12193(eclk, ereset, n_2229_v,(n_165_v|n_872_v), 1'b1,1'b0, n_859_v);
  spice_mux_2 mux_12194(eclk, ereset, n_1209_v,v(n_140_v), 1'b1,1'b0, m2_v);
  spice_mux_2 mux_12195(eclk, ereset, n_1451_v,n_1442_v, 1'b1,1'b0, n_607_v);
  spice_mux_3 mux_12196(eclk, ereset, n_1936_v,n_1914_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_2116_v), n_1968_v);
  spice_mux_3 mux_12197(eclk, ereset, n_858_v,n_851_v,n_1798_v, 1'b1,1'b0,v(n_863_v), n_3452_v);
  spice_mux_3 mux_12198(eclk, ereset, n_853_v,n_2185_v,n_678_v, 1'b1,1'b0,v(n_864_v), n_3453_v);
  spice_mux_2 mux_12199(eclk, ereset, n_1736_v,(n_651_v|n_685_v), 1'b1,1'b0, n_1785_v);
  spice_mux_2 mux_12200(eclk, ereset, n_1961_v,n_724_v, 1'b1,1'b0, n_735_v);
  spice_mux_2 mux_12201(eclk, ereset, n_1579_v,(v(clk_v)|n_543_v), 1'b1,1'b0, n_575_v);
  spice_mux_3 mux_12202(eclk, ereset, n_2556_v,n_2566_v,n_552_v, 1'b1,1'b0,v(n_951_v), n_3547_v);
  spice_mux_2 mux_12203(eclk, ereset, n_2568_v,(n_930_v|n_165_v), 1'b1,1'b0, n_978_v);
  spice_mux_2 mux_12204(eclk, ereset, n_1962_v,n_1789_v, 1'b1,1'b0, n_757_v);
  spice_mux_2 mux_12205(eclk, ereset, n_2560_v,n_2531_v, 1'b1,1'b0, n_2496_v);
  spice_mux_3 mux_12206(eclk, ereset, n_2564_v,n_2557_v,n_553_v, 1'b1,1'b0,v(n_951_v), n_3551_v);
  spice_mux_2 mux_12207(eclk, ereset, n_1119_v,n_1140_v, 1'b1,1'b0, n_131_v);
  spice_mux_2 mux_12208(eclk, ereset, n_1064_v,v(n_84_v), 1'b1,1'b0, n_1037_v);
  spice_mux_2 mux_12209(eclk, ereset, n_1471_v,n_1440_v, 1'b1,1'b0, n_1462_v);
  spice_mux_2 mux_12210(eclk, ereset, n_1964_v,(n_1861_v|v(clk_v)), 1'b1,1'b0, n_740_v);
  spice_mux_3 mux_12211(eclk, ereset, n_742_v,n_743_v,n_1798_v, 1'b1,1'b0,v(n_749_v), n_3396_v);
  spice_mux_2 mux_12212(eclk, ereset, n_1737_v,n_393_v, 1'b1,1'b0, n_680_v);
  spice_mux_3 mux_12213(eclk, ereset, n_1935_v,n_741_v,n_678_v, 1'b1,1'b0,v(n_745_v), n_3395_v);
  spice_mux_2 mux_12214(eclk, ereset, n_1130_v,(n_1147_v|v(clk_v)), 1'b1,1'b0, n_111_v);
  spice_mux_2 mux_12215(eclk, ereset, n_1194_v,v(n_1170_v), 1'b1,1'b0, _t5_v);
  spice_mux_2 mux_12216(eclk, ereset, n_1593_v,n_1602_v, 1'b1,1'b0, n_651_v);
  spice_mux_2 mux_12217(eclk, ereset, n_1766_v,n_1710_v, 1'b1,1'b0, n_643_v);
  spice_mux_3 mux_12218(eclk, ereset, n_977_v,n_976_v,n_1798_v, 1'b1,1'b0,v(n_974_v), n_3549_v);
  spice_mux_2 mux_12219(eclk, ereset, n_2565_v,v(n_956_v), 1'b1,1'b0, n_817_v);
  spice_mux_2 mux_12220(eclk, ereset, n_1292_v,(n_215_v|n_95_v), 1'b1,1'b0, n_110_v);
  spice_mux_3 mux_12221(eclk, ereset, n_975_v,n_2590_v,n_652_v, 1'b1,1'b0,v(n_973_v), n_3550_v);
  spice_mux_2 mux_12222(eclk, ereset, n_1097_v,n_1089_v, 1'b1,1'b0, n_93_v);
  spice_mux_2 mux_12223(eclk, ereset, n_1473_v,n_425_v, 1'b1,1'b0, n_232_v);
  spice_mux_2 mux_12224(eclk, ereset, n_1769_v,n_1764_v, 1'b1,1'b0, n_646_v);
  spice_mux_2 mux_12225(eclk, ereset, n_1335_v,(n_1326_v|v(clk_v)), 1'b1,1'b0, n_162_v);
  spice_mux_2 mux_12226(eclk, ereset, n_1191_v,v(n_89_v), 1'b1,1'b0, _t6_v);
  spice_mux_3 mux_12227(eclk, ereset, n_832_v,v(clk_v),n_604_v, 1'b1,n_2566_v,v(n_951_v), n_968_v);
  spice_mux_2 mux_12228(eclk, ereset, n_2571_v,n_967_v, 1'b1,1'b0, n_943_v);
  spice_mux_2 mux_12229(eclk, ereset, n_1093_v,n_104_v, 1'b1,1'b0, n_105_v);
  spice_mux_2 mux_12230(eclk, ereset, n_1094_v,n_104_v, 1'b1,1'b0, n_66_v);
  spice_mux_3 mux_12231(eclk, ereset, n_2591_v,n_2572_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_1017_v), n_1003_v);
  spice_mux_2 mux_12232(eclk, ereset, n_1103_v,v(n_1076_v), 1'b1,1'b0, n_1040_v);
  spice_mux_2 mux_12233(eclk, ereset, n_1223_v,v(n_1220_v), 1'b1,1'b0, n_165_v);
  spice_mux_3 mux_12234(eclk, ereset, n_976_v,n_977_v,n_1798_v, 1'b1,1'b0,v(n_982_v), n_3554_v);
  spice_mux_3 mux_12235(eclk, ereset, n_2590_v,n_975_v,n_652_v, 1'b1,1'b0,v(n_980_v), n_3553_v);
  spice_mux_2 mux_12236(eclk, ereset, n_1068_v,n_1073_v, 1'b1,1'b0, n_80_v);
  spice_mux_2 mux_12237(eclk, ereset, n_1226_v,(n_170_v|n_165_v), 1'b1,1'b0, n_1207_v);
  spice_mux_2 mux_12238(eclk, ereset, n_1779_v,(n_627_v|n_1774_v), 1'b1,1'b0, n_641_v);
  spice_mux_2 mux_12239(eclk, ereset, n_1969_v,(n_627_v|n_1910_v), 1'b1,1'b0, n_1966_v);
  spice_mux_3 mux_12240(eclk, ereset, n_877_v,n_874_v,n_1798_v, 1'b1,1'b0,v(n_871_v), n_3463_v);
  spice_mux_2 mux_12241(eclk, ereset, n_875_v,(n_825_v|n_855_v), 1'b1,1'b0, n_878_v);
  spice_mux_2 mux_12242(eclk, ereset, n_1788_v,n_573_v, 1'b1,1'b0, n_693_v);
  spice_mux_3 mux_12243(eclk, ereset, n_873_v,n_2250_v,n_652_v, 1'b1,1'b0,v(n_870_v), n_3464_v);
  spice_mux_3 mux_12244(eclk, ereset, n_2224_v,n_2255_v,n_574_v, 1'b1,1'b0,v(n_852_v), n_3467_v);
  spice_mux_2 mux_12245(eclk, ereset, n_1038_v,n_1037_v, 1'b1,1'b0, _iorq_v);
  spice_mux_2 mux_12246(eclk, ereset, n_1599_v,n_520_v, 1'b1,1'b0, n_194_v);
  spice_mux_2 mux_12247(eclk, ereset, n_2636_v,(n_627_v|v(n_2617_v)), 1'b1,1'b0, n_2616_v);
  spice_mux_2 mux_12248(eclk, ereset, n_2616_v,n_2569_v, 1'b1,1'b0, ab4_v);
  spice_mux_3 mux_12249(eclk, ereset, n_760_v,n_771_v,n_1798_v, 1'b1,1'b0,v(n_752_v), n_3399_v);
  spice_mux_3 mux_12250(eclk, ereset, n_987_v,n_996_v,n_1798_v, 1'b1,1'b0,v(n_984_v), n_3558_v);
  spice_mux_3 mux_12251(eclk, ereset, n_95_v,v(clk_v),(n_200_v&n_204_v), 1'b1,n_1262_v,n_1296_v, n_1242_v);
  spice_mux_2 mux_12252(eclk, ereset, n_1790_v,(v(clk_v)|n_649_v), 1'b1,1'b0, n_684_v);
  spice_mux_2 mux_12253(eclk, ereset, n_1301_v,n_1282_v, 1'b1,1'b0, n_222_v);
  spice_mux_3 mux_12254(eclk, ereset, n_2226_v,n_2256_v,n_552_v, 1'b1,1'b0,v(n_852_v), n_3469_v);
  spice_mux_2 mux_12255(eclk, ereset, n_679_v,(v(clk_v)|n_606_v), 1'b1,1'b0, n_678_v);
  spice_mux_2 mux_12256(eclk, ereset, n_1786_v,n_1696_v, 1'b1,1'b0, n_692_v);
  spice_mux_2 mux_12257(eclk, ereset, n_2230_v,n_2223_v, 1'b1,1'b0, n_2186_v);
  spice_mux_2 mux_12258(eclk, ereset, n_1607_v,n_1592_v, 1'b1,1'b0, n_590_v);
  spice_mux_2 mux_12259(eclk, ereset, n_2613_v,(n_978_v|n_165_v), 1'b1,1'b0, n_2615_v);
  spice_mux_3 mux_12260(eclk, ereset, n_2637_v,n_990_v,n_652_v, 1'b1,1'b0,v(n_985_v), n_3560_v);
  spice_mux_2 mux_12261(eclk, ereset, n_653_v,(v(clk_v)|n_620_v), 1'b1,1'b0, n_652_v);
  spice_mux_2 mux_12262(eclk, ereset, n_1620_v,n_1595_v, 1'b1,1'b0, n_574_v);
  spice_mux_3 mux_12263(eclk, ereset, n_2251_v,n_2225_v,(n_393_v&v(clk_v)), 1'b1,1'b0,v(n_2702_v), n_2279_v);
  spice_mux_3 mux_12264(eclk, ereset, n_2227_v,n_866_v,n_553_v, 1'b1,1'b0,v(n_852_v), n_3471_v);
  spice_mux_3 mux_12265(eclk, ereset, n_1991_v,n_761_v,n_678_v, 1'b1,1'b0,v(n_753_v), n_3401_v);
  spice_mux_3 mux_12266(eclk, ereset, n_2663_v,n_2638_v,n_553_v, 1'b1,1'b0,v(n_983_v), n_3557_v);
  spice_mux_3 mux_12267(eclk, ereset, n_2662_v,n_2667_v,n_552_v, 1'b1,1'b0,v(n_983_v), n_3562_v);
  spice_mux_3 mux_12268(eclk, ereset, n_2664_v,n_2668_v,n_646_v, 1'b1,1'b0,v(n_983_v), n_2658_v);
  spice_mux_3 mux_12269(eclk, ereset, n_1990_v,n_1992_v,(v(clk_v)&n_393_v), 1'b1,1'b0,v(n_2320_v), n_1970_v);
  spice_mux_3 mux_12270(eclk, ereset, n_1989_v,n_642_v,(n_2090_v&n_643_v), 1'b1,1'b0,v(n_837_v), n_3404_v);
  spice_mux_2 mux_12271(eclk, ereset, n_1617_v,n_1603_v, 1'b1,1'b0, n_618_v);
  spice_mux_3 mux_12272(eclk, ereset, n_2639_v,n_2660_v,(v(clk_v)&n_393_v), 1'b1,1'b0,v(n_1018_v), n_1004_v);
  spice_mux_2 mux_12273(eclk, ereset, n_1392_v,n_396_v, 1'b1,1'b0, n_65_v);
  spice_mux_3 mux_12274(eclk, ereset, n_874_v,n_877_v,n_1798_v, 1'b1,1'b0,v(n_884_v), n_3473_v);
  spice_mux_3 mux_12275(eclk, ereset, n_2673_v,n_2666_v,n_574_v, 1'b1,1'b0,v(n_983_v), n_3564_v);
  spice_mux_3 mux_12276(eclk, ereset, n_2250_v,n_873_v,n_652_v, 1'b1,1'b0,v(n_880_v), n_3472_v);
  spice_mux_3 mux_12277(eclk, ereset, n_996_v,n_987_v,n_1798_v, 1'b1,1'b0,v(n_998_v), n_3569_v);
  spice_mux_3 mux_12278(eclk, ereset, n_990_v,n_2637_v,n_652_v, 1'b1,1'b0,v(n_999_v), n_3570_v);
  spice_mux_3 mux_12279(eclk, ereset, n_832_v,v(clk_v),n_604_v, 1'b1,n_2256_v,v(n_852_v), n_868_v);
  spice_mux_2 mux_12280(eclk, ereset, n_2273_v,n_869_v, 1'b1,1'b0, n_844_v);
  spice_mux_2 mux_12281(eclk, ereset, n_1625_v,n_1587_v, 1'b1,1'b0, n_552_v);
  spice_mux_2 mux_12282(eclk, ereset, n_655_v,(v(clk_v)|n_599_v), 1'b1,1'b0, n_654_v);
  spice_mux_3 mux_12283(eclk, ereset, n_95_v,n_204_v,v(clk_v), 1'b1,n_200_v,n_1267_v, n_1243_v);
  spice_mux_2 mux_12284(eclk, ereset, n_397_v,n_1394_v, 1'b1,1'b0, n_1393_v);
  spice_mux_2 mux_12285(eclk, ereset, n_656_v,(v(clk_v)|n_602_v), 1'b1,1'b0, n_657_v);
  spice_mux_2 mux_12286(eclk, ereset, n_659_v,(v(clk_v)|n_1738_v), 1'b1,1'b0, n_658_v);
  spice_mux_3 mux_12287(eclk, ereset, n_95_v,n_204_v,v(clk_v), 1'b1,n_1248_v,n_1273_v, n_1245_v);
  spice_mux_2 mux_12288(eclk, ereset, n_1338_v,(n_250_v|n_165_v), 1'b1,1'b0, n_1336_v);
  spice_mux_2 mux_12289(eclk, ereset, n_660_v,(v(clk_v)|n_1739_v), 1'b1,1'b0, n_661_v);
  spice_mux_2 mux_12290(eclk, ereset, n_663_v,(v(clk_v)|n_1740_v), 1'b1,1'b0, n_662_v);
  spice_mux_2 mux_12291(eclk, ereset, n_1482_v,n_1469_v, 1'b1,1'b0, n_479_v);
  spice_mux_2 mux_12292(eclk, ereset, n_1340_v,(v(n_244_v)|n_255_v), 1'b1,1'b0, n_326_v);
  spice_mux_2 mux_12293(eclk, ereset, n_664_v,(v(clk_v)|n_1741_v), 1'b1,1'b0, n_665_v);
  spice_mux_3 mux_12294(eclk, ereset, n_771_v,n_760_v,n_1798_v, 1'b1,1'b0,v(n_774_v), n_3405_v);
  spice_mux_3 mux_12295(eclk, ereset, n_761_v,n_1991_v,n_678_v, 1'b1,1'b0,v(n_775_v), n_3406_v);
  spice_mux_2 mux_12296(eclk, ereset, n_667_v,(v(clk_v)|n_1742_v), 1'b1,1'b0, n_666_v);
  spice_mux_2 mux_12297(eclk, ereset, n_1344_v,v(n_259_v), 1'b1,1'b0, m1_v);
  spice_mux_2 mux_12298(eclk, ereset, n_1631_v,n_1600_v, 1'b1,1'b0, n_553_v);
  spice_mux_3 mux_12299(eclk, ereset, n_888_v,n_895_v,n_1798_v, 1'b1,1'b0,v(n_885_v), n_3477_v);
  spice_mux_2 mux_12300(eclk, ereset, n_668_v,(v(clk_v)|n_1743_v), 1'b1,1'b0, n_669_v);
  spice_mux_2 mux_12301(eclk, ereset, n_671_v,(v(clk_v)|n_1744_v), 1'b1,1'b0, n_670_v);
  spice_mux_2 mux_12302(eclk, ereset, n_1401_v,n_371_v, 1'b1,1'b0, n_1385_v);
  spice_mux_2 mux_12303(eclk, ereset, n_1149_v,n_1111_v, 1'b1,1'b0, n_129_v);
  spice_mux_2 mux_12304(eclk, ereset, n_672_v,(v(clk_v)|n_1745_v), 1'b1,1'b0, n_673_v);
  spice_mux_2 mux_12305(eclk, ereset, n_675_v,(v(clk_v)|n_1746_v), 1'b1,1'b0, n_674_v);
  spice_mux_2 mux_12306(eclk, ereset, n_1638_v,n_1598_v, 1'b1,1'b0, n_612_v);
  spice_mux_2 mux_12307(eclk, ereset, n_1627_v,n_1532_v, 1'b1,1'b0, n_558_v);
  spice_mux_2 mux_12308(eclk, ereset, n_676_v,(v(clk_v)|n_1747_v), 1'b1,1'b0, n_677_v);
  spice_mux_2 mux_12309(eclk, ereset, n_1339_v,v(n_240_v), 1'b1,1'b0, n_327_v);
  spice_mux_2 mux_12310(eclk, ereset, n_1008_v,(n_825_v|n_997_v), 1'b1,1'b0, n_827_v);
  spice_mux_3 mux_12311(eclk, ereset, n_2680_v,n_2690_v,n_574_v, 1'b1,1'b0,v(n_995_v), n_3581_v);
  spice_mux_2 mux_12312(eclk, ereset, n_1070_v,(n_113_v|(n_79_v&n_122_v)), 1'b1,1'b0, n_78_v);
  spice_mux_2 mux_12313(eclk, ereset, n_1492_v,n_1472_v, 1'b1,1'b0, n_548_v);
  spice_mux_3 mux_12314(eclk, ereset, n_2677_v,n_2679_v,n_87_v, 1'b1,1'b0,v(n_485_v), n_3579_v);
  spice_mux_2 mux_12315(eclk, ereset, n_1634_v,n_1565_v, 1'b1,1'b0, n_551_v);
  spice_mux_3 mux_12316(eclk, ereset, n_2682_v,n_2691_v,n_552_v, 1'b1,1'b0,v(n_995_v), n_3583_v);
  spice_mux_3 mux_12317(eclk, ereset, n_2300_v,n_890_v,n_652_v, 1'b1,1'b0,v(n_886_v), n_3479_v);
  spice_mux_2 mux_12318(eclk, ereset, n_2683_v,n_2678_v, 1'b1,1'b0, n_2659_v);
  spice_mux_3 mux_12319(eclk, ereset, n_2299_v,n_2301_v,(v(clk_v)&n_393_v), 1'b1,1'b0,v(n_2703_v), n_2280_v);
  spice_mux_2 mux_12320(eclk, ereset, n_1626_v,v(n_1586_v), 1'b1,1'b0, n_549_v);
  spice_mux_3 mux_12321(eclk, ereset, n_2687_v,n_2681_v,n_553_v, 1'b1,1'b0,v(n_995_v), n_3584_v);
  spice_mux_2 mux_12322(eclk, ereset, n_2688_v,v(n_1001_v), 1'b1,1'b0, n_830_v);
  spice_mux_2 mux_12323(eclk, ereset, n_2014_v,(n_778_v|n_627_v), 1'b1,1'b0, n_2044_v);
  spice_mux_2 mux_12324(eclk, ereset, n_1400_v,n_326_v, 1'b1,1'b0, n_1354_v);
  spice_mux_3 mux_12325(eclk, ereset, n_832_v,v(clk_v),n_604_v, 1'b1,n_2691_v,v(n_995_v), n_1007_v);
  spice_mux_2 mux_12326(eclk, ereset, n_2693_v,n_1006_v, 1'b1,1'b0, n_989_v);
  spice_mux_2 mux_12327(eclk, ereset, n_2696_v,(v(n_1009_v)|n_627_v), 1'b1,1'b0, n_2695_v);
  spice_mux_2 mux_12328(eclk, ereset, n_1303_v,n_1259_v, 1'b1,1'b0, n_265_v);
  spice_mux_2 mux_12329(eclk, ereset, n_2699_v,v(n_486_v), 1'b1,1'b0, n_883_v);
  spice_mux_2 mux_12330(eclk, ereset, n_2697_v,(n_1011_v|n_165_v), 1'b1,1'b0, n_2706_v);
  spice_mux_2 mux_12331(eclk, ereset, v(ex_bcdehl_v),v(n_1773_v), 1'b1,1'b0, n_634_v);
  spice_mux_2 mux_12332(eclk, ereset, n_2707_v,(n_165_v|n_1000_v), 1'b1,1'b0, n_1011_v);
  spice_mux_2 mux_12333(eclk, ereset, n_2708_v,(n_1026_v|n_627_v), 1'b1,1'b0, n_2741_v);
  spice_mux_2 mux_12334(eclk, ereset, n_1197_v,v(n_147_v), 1'b1,1'b0, _t2_v);
  spice_mux_2 mux_12335(eclk, ereset, n_1803_v,(v(clk_v)|n_589_v), 1'b1,1'b0, n_695_v);
  spice_mux_2 mux_12336(eclk, ereset, n_1236_v,v(n_1228_v), 1'b1,1'b0, m3_v);
  spice_mux_2 mux_12337(eclk, ereset, n_1348_v,n_357_v, 1'b1,1'b0, n_1347_v);
  spice_mux_3 mux_12338(eclk, ereset, n_895_v,n_888_v,n_1798_v, 1'b1,1'b0,v(n_901_v), n_3484_v);
  spice_mux_2 mux_12339(eclk, ereset, n_1795_v,(v(clk_v)|n_588_v), 1'b1,1'b0, n_1798_v);
  spice_mux_2 mux_12340(eclk, ereset, n_1796_v,(v(clk_v)|n_590_v), 1'b1,1'b0, n_1799_v);
  spice_mux_3 mux_12341(eclk, ereset, n_890_v,n_2300_v,n_652_v, 1'b1,1'b0,v(n_902_v), n_3486_v);
  spice_mux_2 mux_12342(eclk, ereset, n_1797_v,(v(clk_v)|n_1674_v), 1'b1,1'b0, n_1800_v);
  spice_mux_3 mux_12343(eclk, ereset, n_2333_v,n_2323_v,n_553_v, 1'b1,1'b0,v(n_889_v), n_3482_v);
  spice_mux_3 mux_12344(eclk, ereset, n_2336_v,n_2324_v,n_87_v, 1'b1,1'b0,v(n_486_v), n_3483_v);
  spice_mux_3 mux_12345(eclk, ereset, n_2332_v,n_2335_v,n_552_v, 1'b1,1'b0,v(n_889_v), n_3485_v);
  spice_mux_3 mux_12346(eclk, ereset, n_2334_v,n_2339_v,n_646_v, 1'b1,1'b0,v(n_889_v), n_2328_v);
  spice_mux_3 mux_12347(eclk, ereset, n_782_v,n_781_v,n_1798_v, 1'b1,1'b0,v(n_777_v), n_3417_v);
  spice_mux_2 mux_12348(eclk, ereset, n_1495_v,n_1468_v, 1'b1,1'b0, n_484_v);
  spice_mux_3 mux_12349(eclk, ereset, n_780_v,n_2036_v,n_678_v, 1'b1,1'b0,v(n_776_v), n_3418_v);
  spice_mux_2 mux_12350(eclk, ereset, n_2725_v,(n_627_v|v(n_2700_v)), 1'b1,1'b0, n_2731_v);
  spice_mux_2 mux_12351(eclk, ereset, n_2726_v,(v(n_2705_v)|n_627_v), 1'b1,1'b0, n_2736_v);
  spice_mux_2 mux_12352(eclk, ereset, n_2727_v,(v(n_2701_v)|n_627_v), 1'b1,1'b0, n_2732_v);
  spice_mux_2 mux_12353(eclk, ereset, n_2728_v,(n_627_v|v(n_2702_v)), 1'b1,1'b0, n_2733_v);
  spice_mux_2 mux_12354(eclk, ereset, n_2729_v,(v(n_2703_v)|n_627_v), 1'b1,1'b0, n_2734_v);
  spice_mux_2 mux_12355(eclk, ereset, n_2730_v,(n_627_v|v(n_2704_v)), 1'b1,1'b0, n_2735_v);
  spice_mux_2 mux_12356(eclk, ereset, n_2017_v,n_610_v, 1'b1,1'b0, n_793_v);
  spice_mux_2 mux_12357(eclk, ereset, v(n_124_v),((v(n_1080_v)|n_1081_v)|(n_1082_v&v(clk_v))), 1'b1,1'b0, n_82_v);
  spice_mux_2 mux_12358(eclk, ereset, n_1293_v,n_224_v, 1'b1,1'b0, n_72_v);
  spice_mux_2 mux_12359(eclk, ereset, n_1402_v,n_381_v, 1'b1,1'b0, n_406_v);
  spice_mux_2 mux_12360(eclk, ereset, n_2719_v,(n_1012_v|n_627_v), 1'b1,1'b0, n_2742_v);
  spice_mux_2 mux_12361(eclk, ereset, n_1289_v,n_1189_v, 1'b1,1'b0, n_270_v);
  spice_mux_2 mux_12362(eclk, ereset, n_1642_v,n_1606_v, 1'b1,1'b0, n_546_v);
  spice_mux_2 mux_12363(eclk, ereset, n_1635_v,n_1577_v, 1'b1,1'b0, n_599_v);
  spice_mux_2 mux_12364(eclk, ereset, n_2709_v,(n_1013_v|n_627_v), 1'b1,1'b0, n_2755_v);
  spice_mux_2 mux_12365(eclk, ereset, n_2710_v,(n_627_v|n_1021_v), 1'b1,1'b0, n_2743_v);
  spice_mux_2 mux_12366(eclk, ereset, n_2711_v,(n_1022_v|n_627_v), 1'b1,1'b0, n_2744_v);
  spice_mux_2 mux_12367(eclk, ereset, n_2712_v,(n_627_v|n_1023_v), 1'b1,1'b0, n_2745_v);
  spice_mux_2 mux_12368(eclk, ereset, n_2713_v,(n_1024_v|n_627_v), 1'b1,1'b0, n_2746_v);
  spice_mux_2 mux_12369(eclk, ereset, n_2714_v,(n_627_v|n_1025_v), 1'b1,1'b0, n_2747_v);
  spice_mux_2 mux_12370(eclk, ereset, n_2749_v,(v(n_1020_v)|n_627_v), 1'b1,1'b0, n_2748_v);
  spice_mux_3 mux_12371(eclk, ereset, n_2342_v,n_2337_v,n_574_v, 1'b1,1'b0,v(n_889_v), n_3487_v);
  spice_mux_2 mux_12372(eclk, ereset, n_2750_v,(n_627_v|v(n_1014_v)), 1'b1,1'b0, n_2756_v);
  spice_mux_2 mux_12373(eclk, ereset, n_2716_v,(n_627_v|n_1015_v), 1'b1,1'b0, n_2757_v);
  spice_mux_2 mux_12374(eclk, ereset, n_2717_v,(n_1016_v|n_627_v), 1'b1,1'b0, n_2758_v);
  spice_mux_2 mux_12375(eclk, ereset, n_2752_v,(v(n_1017_v)|n_627_v), 1'b1,1'b0, n_2751_v);
  spice_mux_2 mux_12376(eclk, ereset, n_357_v,n_1348_v, 1'b1,1'b0, n_374_v);
  spice_mux_2 mux_12377(eclk, ereset, n_2753_v,(n_627_v|v(n_1018_v)), 1'b1,1'b0, n_2754_v);
  spice_mux_2 mux_12378(eclk, ereset, n_2718_v,(n_627_v|n_1019_v), 1'b1,1'b0, n_2759_v);
  spice_mux_2 mux_12379(eclk, ereset, n_1497_v,n_1467_v, 1'b1,1'b0, n_330_v);
  spice_mux_2 mux_12380(eclk, ereset, n_2695_v,n_2741_v, 1'b1,1'b0, ab5_v);
  spice_mux_2 mux_12381(eclk, ereset, n_2731_v,n_2742_v, 1'b1,1'b0, ab6_v);
  spice_mux_2 mux_12382(eclk, ereset, n_2732_v,n_2743_v, 1'b1,1'b0, ab7_v);
  spice_mux_2 mux_12383(eclk, ereset, n_2733_v,n_2744_v, 1'b1,1'b0, ab8_v);
  spice_mux_2 mux_12384(eclk, ereset, n_2734_v,n_2745_v, 1'b1,1'b0, ab9_v);
  spice_mux_2 mux_12385(eclk, ereset, n_2735_v,n_2746_v, 1'b1,1'b0, ab10_v);
  spice_mux_2 mux_12386(eclk, ereset, n_2736_v,n_2747_v, 1'b1,1'b0, ab11_v);
  spice_mux_2 mux_12387(eclk, ereset, n_2748_v,n_2755_v, 1'b1,1'b0, ab12_v);
  spice_mux_2 mux_12388(eclk, ereset, n_2756_v,n_2757_v, 1'b1,1'b0, ab13_v);
  spice_mux_2 mux_12389(eclk, ereset, n_2751_v,n_2758_v, 1'b1,1'b0, ab14_v);
  spice_mux_2 mux_12390(eclk, ereset, n_2754_v,n_2759_v, 1'b1,1'b0, ab15_v);
  spice_mux_2 mux_12391(eclk, ereset, n_1403_v,n_420_v, 1'b1,1'b0, n_387_v);
  spice_mux_3 mux_12392(eclk, ereset, n_476_v,n_474_v,n_474_v, 1'b0,v(n_475_v),v(n_475_v), n_474_v);
  spice_mux_3 mux_12393(eclk, ereset, n_474_v,n_1491_v,n_1491_v, 1'b0,v(n_475_v),v(n_475_v), n_1491_v);
  spice_mux_3 mux_12394(eclk, ereset, n_471_v,n_471_v,n_476_v, 1'b0,n_476_v,v(n_475_v), n_3014_v);
  spice_mux_3 mux_12395(eclk, ereset, n_474_v,n_1501_v,n_1501_v, 1'b0,v(n_475_v),v(n_475_v), n_1501_v);
  spice_mux_2 mux_12396(eclk, ereset, n_476_v,n_476_v, v(n_475_v),v(n_475_v), n_476_v);
  spice_mux_3 mux_12397(eclk, ereset, v(clk_v),n_207_v,(n_188_v|n_95_v), n_1239_v,v(n_248_v),1'b0, n_206_v);
  spice_mux_3 mux_12398(eclk, ereset, n_95_v,v(clk_v),n_180_v, 1'b0,n_1268_v,v(n_248_v), n_205_v);
  spice_mux_3 mux_12399(eclk, ereset, n_1196_v,n_82_v,n_133_v, n_1181_v,n_1150_v,v(n_138_v), n_123_v);
  spice_mux_3 mux_12400(eclk, ereset, n_133_v,n_1308_v,n_82_v, v(n_196_v),n_1288_v,n_1257_v, n_195_v);
  spice_mux_2 mux_12401(eclk, ereset, n_521_v,v(clk_v), n_1645_v,n_1640_v, n_1615_v);
  spice_mux_2 mux_12402(eclk, ereset, v(clk_v),n_611_v, n_1637_v,n_688_v, n_1682_v);
  spice_mux_2 mux_12403(eclk, ereset, ex_dehl_combined_v,n_1713_v, n_601_v,v(n_616_v), n_1705_v);
  spice_mux_2 mux_12404(eclk, ereset, n_1708_v,ex_dehl_combined_v, n_601_v,v(n_616_v), n_1706_v);
  spice_mux_3 mux_12405(eclk, ereset, n_95_v,v(clk_v),n_204_v, 1'b0,n_1182_v,n_130_v, n_1145_v);
  spice_mux_2 mux_12406(eclk, ereset, n_695_v,v(clk_v), n_1828_v,n_1856_v, n_1830_v);
  spice_mux_2 mux_12407(eclk, ereset, n_1354_v,n_326_v, v(n_138_v),n_357_v, n_1350_v);
  spice_mux_3 mux_12408(eclk, ereset, n_575_v,n_712_v,v(clk_v), v(n_525_v),n_1944_v,n_1959_v, n_729_v);
  spice_mux_2 mux_12409(eclk, ereset, v(clk_v),n_695_v, n_1887_v,n_1906_v, n_1909_v);
  spice_mux_2 mux_12410(eclk, ereset, n_326_v,n_1354_v, n_373_v,v(n_196_v), n_1360_v);
  spice_mux_2 mux_12411(eclk, ereset, n_695_v,v(clk_v), n_1929_v,n_1963_v, n_1931_v);
  spice_mux_3 mux_12412(eclk, ereset, n_82_v,n_2016_v,n_133_v, n_2015_v,n_788_v,v(n_380_v), n_751_v);
  spice_mux_3 mux_12413(eclk, ereset, n_82_v,n_1367_v,n_133_v, n_1349_v,n_1362_v,v(n_370_v), n_358_v);
  spice_mux_2 mux_12414(eclk, ereset, n_1354_v,n_326_v, v(n_412_v),n_376_v, n_1366_v);
  spice_mux_2 mux_12415(eclk, ereset, v(clk_v),n_695_v, n_1993_v,n_2012_v, n_2013_v);
  spice_mux_2 mux_12416(eclk, ereset, n_695_v,v(clk_v), n_2033_v,n_2060_v, n_2034_v);
  spice_mux_2 mux_12417(eclk, ereset, n_1354_v,n_326_v, v(n_380_v),n_379_v, n_1370_v);
  spice_mux_2 mux_12418(eclk, ereset, v(clk_v),n_695_v, n_2089_v,n_2113_v, n_2114_v);
  spice_mux_2 mux_12419(eclk, ereset, n_695_v,v(clk_v), n_2133_v,n_2157_v, n_2134_v);
  spice_mux_2 mux_12420(eclk, ereset, v(clk_v),n_695_v, n_2190_v,n_2221_v, n_2222_v);
  spice_mux_2 mux_12421(eclk, ereset, n_1354_v,n_326_v, v(n_370_v),n_382_v, n_1375_v);
  spice_mux_2 mux_12422(eclk, ereset, n_831_v,n_747_v, n_2191_v,v(n_2211_v), n_865_v);
  spice_mux_3 mux_12423(eclk, ereset, n_2389_v,n_82_v,n_133_v, n_2336_v,n_2277_v,v(n_486_v), n_872_v);
  spice_mux_2 mux_12424(eclk, ereset, n_695_v,v(clk_v), n_2246_v,n_2275_v, n_2248_v);
  spice_mux_2 mux_12425(eclk, ereset, n_1354_v,n_326_v, v(n_480_v),n_388_v, n_1380_v);
  spice_mux_2 mux_12426(eclk, ereset, n_695_v,v(clk_v), n_2325_v,n_2303_v, n_2329_v);
  spice_mux_2 mux_12427(eclk, ereset, n_1354_v,n_326_v, v(n_485_v),n_392_v, n_1388_v);
  spice_mux_2 mux_12428(eclk, ereset, n_695_v,v(clk_v), n_2359_v,n_2387_v, n_2361_v);
  spice_mux_2 mux_12429(eclk, ereset, n_831_v,n_747_v, n_2334_v,v(n_2338_v), n_912_v);
  spice_mux_2 mux_12430(eclk, ereset, n_1354_v,n_326_v, v(n_486_v),n_397_v, n_1395_v);
  spice_mux_2 mux_12431(eclk, ereset, v(clk_v),n_695_v, n_2424_v,n_2446_v, n_2448_v);
  spice_mux_3 mux_12432(eclk, ereset, n_2425_v,n_133_v,n_82_v, n_2445_v,v(n_480_v),n_2535_v, n_930_v);
  spice_mux_2 mux_12433(eclk, ereset, n_695_v,v(clk_v), n_2464_v,n_2495_v, n_2465_v);
  spice_mux_2 mux_12434(eclk, ereset, n_831_v,n_747_v, n_2500_v,v(n_2504_v), n_960_v);
  spice_mux_2 mux_12435(eclk, ereset, v(clk_v),n_695_v, n_2536_v,n_2559_v, n_2562_v);
  spice_mux_2 mux_12436(eclk, ereset, n_695_v,v(clk_v), n_2587_v,n_2612_v, n_2588_v);
  spice_mux_3 mux_12437(eclk, ereset, n_133_v,n_82_v,n_1407_v, v(n_412_v),n_1422_v,n_1408_v, n_414_v);
  spice_mux_2 mux_12438(eclk, ereset, v(clk_v),n_695_v, n_2640_v,n_2671_v, n_2674_v);
  spice_mux_2 mux_12439(eclk, ereset, n_831_v,n_747_v, n_2664_v,v(n_816_v), n_1002_v);
  spice_mux_3 mux_12440(eclk, ereset, n_2669_v,n_133_v,n_82_v, n_2677_v,v(n_485_v),n_1010_v, n_1000_v);
  spice_mux_2 mux_12441(eclk, ereset, n_95_v,v(clk_v), 1'b0,n_1215_v, n_179_v);
  spice_mux_3 mux_12442(eclk, ereset, n_1460_v,n_712_v,n_1805_v, n_683_v,v(n_647_v),v(n_700_v), n_3358_v);
  spice_mux_3 mux_12443(eclk, ereset, n_1930_v,n_735_v,n_643_v, v(n_726_v),v(n_545_v),v(n_525_v), n_1942_v);

  spice_node_4 n_n_779(eclk, ereset, n_779_port_3,n_779_port_4,n_779_port_5,n_779_port_8, n_779_v);
  spice_node_4 n_n_791(eclk, ereset, n_791_port_0,n_791_port_1,n_791_port_3,n_791_port_4, n_791_v);
  spice_node_2 n_n_1498(eclk, ereset, n_1498_port_2,n_1498_port_3, n_1498_v);
  spice_node_4 n_n_703(eclk, ereset, n_703_port_0,n_703_port_3,n_703_port_4,n_703_port_5, n_703_v);
  spice_node_4 n_n_907(eclk, ereset, n_907_port_0,n_907_port_3,n_907_port_4,n_907_port_5, n_907_v);
  spice_node_3 n_db0(eclk, ereset, db0_port_0,db0_port_1,db0_port_3, db0_v);
  spice_node_3 n_db7(eclk, ereset, db7_port_0,db7_port_2,db7_port_3, db7_v);
  spice_node_6 n_n_783(eclk, ereset, n_783_port_5,n_783_port_6,n_783_port_7,n_783_port_8,n_783_port_9,n_783_port_10, n_783_v);
  spice_node_3 n_db1(eclk, ereset, db1_port_0,db1_port_2,db1_port_3, db1_v);
  spice_node_2 n_n_380(eclk, ereset, n_380_port_0,n_380_port_2, n_380_v);
  spice_node_2 n_n_480(eclk, ereset, n_480_port_0,n_480_port_7, n_480_v);
  spice_node_2 n_n_485(eclk, ereset, n_485_port_0,n_485_port_7, n_485_v);
  spice_node_2 n_n_486(eclk, ereset, n_486_port_0,n_486_port_6, n_486_v);
  spice_node_4 n_n_713(eclk, ereset, n_713_port_0,n_713_port_1,n_713_port_3,n_713_port_4, n_713_v);
  spice_node_6 n_n_545(eclk, ereset, n_545_port_4,n_545_port_8,n_545_port_10,n_545_port_11,n_545_port_12,n_545_port_14, n_545_v);
  spice_node_4 n_n_917(eclk, ereset, n_917_port_0,n_917_port_1,n_917_port_3,n_917_port_4, n_917_v);
  spice_node_4 n_n_798(eclk, ereset, n_798_port_0,n_798_port_2,n_798_port_3,n_798_port_4, n_798_v);
  spice_node_2 n_n_370(eclk, ereset, n_370_port_0,n_370_port_4, n_370_v);
  spice_node_2 n_n_196(eclk, ereset, n_196_port_0,n_196_port_4, n_196_v);
  spice_node_2 n_n_412(eclk, ereset, n_412_port_0,n_412_port_4, n_412_v);
  spice_node_2 n_n_138(eclk, ereset, n_138_port_0,n_138_port_3, n_138_v);
  spice_node_4 n_n_790(eclk, ereset, n_790_port_0,n_790_port_1,n_790_port_3,n_790_port_5, n_790_v);
  spice_node_4 n_n_922(eclk, ereset, n_922_port_0,n_922_port_2,n_922_port_3,n_922_port_4, n_922_v);
  spice_node_4 n_n_806(eclk, ereset, n_806_port_0,n_806_port_3,n_806_port_4,n_806_port_5, n_806_v);
  spice_node_7 n_n_525(eclk, ereset, n_525_port_3,n_525_port_7,n_525_port_8,n_525_port_9,n_525_port_11,n_525_port_13,n_525_port_15, n_525_v);
  spice_node_6 n_n_808(eclk, ereset, n_808_port_5,n_808_port_6,n_808_port_7,n_808_port_8,n_808_port_9,n_808_port_10, n_808_v);
  spice_node_3 n_n_2338(eclk, ereset, n_2338_port_0,n_2338_port_3,n_2338_port_5, n_2338_v);
  spice_node_6 n_n_796(eclk, ereset, n_796_port_5,n_796_port_6,n_796_port_7,n_796_port_8,n_796_port_9,n_796_port_10, n_796_v);
  spice_node_4 n_n_933(eclk, ereset, n_933_port_0,n_933_port_3,n_933_port_4,n_933_port_5, n_933_v);
  spice_node_4 n_n_714(eclk, ereset, n_714_port_0,n_714_port_2,n_714_port_3,n_714_port_4, n_714_v);
  spice_node_3 n_db6(eclk, ereset, db6_port_0,db6_port_1,db6_port_3, db6_v);
  spice_node_3 n_n_248(eclk, ereset, n_248_port_0,n_248_port_25,n_248_port_26, n_248_v);
  spice_node_2 n_n_1332(eclk, ereset, n_1332_port_1,n_1332_port_2, n_1332_v);
  spice_node_2 n_n_73(eclk, ereset, n_73_port_4,n_73_port_6, n_73_v);
  spice_node_5 n_n_528(eclk, ereset, n_528_port_0,n_528_port_1,n_528_port_3,n_528_port_6,n_528_port_7, n_528_v);
  spice_node_4 n_n_810(eclk, ereset, n_810_port_0,n_810_port_3,n_810_port_4,n_810_port_5, n_810_v);
  spice_node_4 n_n_936(eclk, ereset, n_936_port_0,n_936_port_3,n_936_port_4,n_936_port_5, n_936_v);
  spice_node_4 n_n_731(eclk, ereset, n_731_port_0,n_731_port_3,n_731_port_4,n_731_port_5, n_731_v);
  spice_node_2 n_n_616(eclk, ereset, n_616_port_0,n_616_port_1, n_616_v);
  spice_node_6 n_n_803(eclk, ereset, n_803_port_5,n_803_port_6,n_803_port_7,n_803_port_8,n_803_port_9,n_803_port_10, n_803_v);
  spice_node_4 n_n_944(eclk, ereset, n_944_port_0,n_944_port_2,n_944_port_3,n_944_port_4, n_944_v);
  spice_node_5 n_n_716(eclk, ereset, n_716_port_0,n_716_port_3,n_716_port_4,n_716_port_7,n_716_port_8, n_716_v);
  spice_node_4 n_n_947(eclk, ereset, n_947_port_0,n_947_port_2,n_947_port_3,n_947_port_4, n_947_v);
  spice_node_4 n_n_953(eclk, ereset, n_953_port_0,n_953_port_1,n_953_port_3,n_953_port_4, n_953_v);
  spice_node_4 n_n_841(eclk, ereset, n_841_port_0,n_841_port_1,n_841_port_3,n_841_port_4, n_841_v);
  spice_node_3 n_db2(eclk, ereset, db2_port_0,db2_port_1,db2_port_3, db2_v);
  spice_node_4 n_n_845(eclk, ereset, n_845_port_0,n_845_port_2,n_845_port_3,n_845_port_4, n_845_v);
  spice_node_4 n_n_958(eclk, ereset, n_958_port_0,n_958_port_2,n_958_port_3,n_958_port_4, n_958_v);
  spice_node_5 n_n_755(eclk, ereset, n_755_port_5,n_755_port_6,n_755_port_7,n_755_port_8,n_755_port_9, n_755_v);
  spice_node_4 n_n_846(eclk, ereset, n_846_port_0,n_846_port_2,n_846_port_3,n_846_port_4, n_846_v);
  spice_node_4 n_n_739(eclk, ereset, n_739_port_0,n_739_port_3,n_739_port_4,n_739_port_5, n_739_v);
  spice_node_4 n_n_850(eclk, ereset, n_850_port_0,n_850_port_2,n_850_port_3,n_850_port_4, n_850_v);
  spice_node_4 n_n_969(eclk, ereset, n_969_port_0,n_969_port_3,n_969_port_4,n_969_port_5, n_969_v);
  spice_node_4 n_n_863(eclk, ereset, n_863_port_0,n_863_port_3,n_863_port_4,n_863_port_5, n_863_v);
  spice_node_3 n_db5(eclk, ereset, db5_port_0,db5_port_1,db5_port_3, db5_v);
  spice_node_5 n_n_526(eclk, ereset, n_526_port_0,n_526_port_3,n_526_port_6,n_526_port_7,n_526_port_8, n_526_v);
  spice_node_3 n_db3(eclk, ereset, db3_port_0,db3_port_2,db3_port_3, db3_v);
  spice_node_4 n_n_749(eclk, ereset, n_749_port_0,n_749_port_1,n_749_port_3,n_749_port_4, n_749_v);
  spice_node_4 n_n_974(eclk, ereset, n_974_port_0,n_974_port_3,n_974_port_4,n_974_port_5, n_974_v);
  spice_node_6 n_n_836(eclk, ereset, n_836_port_5,n_836_port_6,n_836_port_7,n_836_port_8,n_836_port_9,n_836_port_10, n_836_v);
  spice_node_3 n_n_2504(eclk, ereset, n_2504_port_0,n_2504_port_3,n_2504_port_5, n_2504_v);
  spice_node_4 n_n_966(eclk, ereset, n_966_port_0,n_966_port_2,n_966_port_3,n_966_port_4, n_966_v);
  spice_node_4 n_n_982(eclk, ereset, n_982_port_0,n_982_port_1,n_982_port_3,n_982_port_4, n_982_v);
  spice_node_5 n_n_681(eclk, ereset, n_681_port_5,n_681_port_6,n_681_port_7,n_681_port_8,n_681_port_9, n_681_v);
  spice_node_4 n_n_871(eclk, ereset, n_871_port_0,n_871_port_3,n_871_port_4,n_871_port_5, n_871_v);
  spice_node_4 n_n_752(eclk, ereset, n_752_port_0,n_752_port_2,n_752_port_3,n_752_port_4, n_752_v);
  spice_node_4 n_n_984(eclk, ereset, n_984_port_0,n_984_port_2,n_984_port_3,n_984_port_4, n_984_v);
  spice_node_0 n_n_562(eclk, ereset,  n_562_v);
  spice_node_4 n_n_993(eclk, ereset, n_993_port_0,n_993_port_2,n_993_port_3,n_993_port_4, n_993_v);
  spice_node_5 n_n_839(eclk, ereset, n_839_port_5,n_839_port_6,n_839_port_7,n_839_port_8,n_839_port_9, n_839_v);
  spice_node_3 n_n_2211(eclk, ereset, n_2211_port_0,n_2211_port_3,n_2211_port_5, n_2211_v);
  spice_node_4 n_n_884(eclk, ereset, n_884_port_0,n_884_port_1,n_884_port_3,n_884_port_4, n_884_v);
  spice_node_4 n_n_998(eclk, ereset, n_998_port_0,n_998_port_3,n_998_port_4,n_998_port_5, n_998_v);
  spice_node_4 n_n_770(eclk, ereset, n_770_port_2,n_770_port_4,n_770_port_5,n_770_port_6, n_770_v);
  spice_node_4 n_n_774(eclk, ereset, n_774_port_0,n_774_port_3,n_774_port_4,n_774_port_5, n_774_v);
  spice_node_4 n_n_885(eclk, ereset, n_885_port_0,n_885_port_2,n_885_port_3,n_885_port_4, n_885_v);
  spice_node_3 n_n_816(eclk, ereset, n_816_port_0,n_816_port_4,n_816_port_6, n_816_v);
  spice_node_4 n_n_1005(eclk, ereset, n_1005_port_3,n_1005_port_4,n_1005_port_5,n_1005_port_6, n_1005_v);
  spice_node_6 n_n_772(eclk, ereset, n_772_port_5,n_772_port_6,n_772_port_7,n_772_port_8,n_772_port_9,n_772_port_10, n_772_v);
  spice_node_1 n_clk(eclk, ereset, clk_port_403, clk_v);
  spice_node_2 n_ex_bcdehl(eclk, ereset, ex_bcdehl_port_5,ex_bcdehl_port_8, ex_bcdehl_v);
  spice_node_4 n_n_897(eclk, ereset, n_897_port_0,n_897_port_2,n_897_port_3,n_897_port_4, n_897_v);
  spice_node_4 n_n_901(eclk, ereset, n_901_port_0,n_901_port_2,n_901_port_3,n_901_port_5, n_901_v);
  spice_node_4 n_n_899(eclk, ereset, n_899_port_0,n_899_port_2,n_899_port_3,n_899_port_4, n_899_v);
  spice_node_5 n_n_697(eclk, ereset, n_697_port_0,n_697_port_1,n_697_port_3,n_697_port_4,n_697_port_5, n_697_v);
  spice_node_4 n_n_777(eclk, ereset, n_777_port_0,n_777_port_3,n_777_port_4,n_777_port_5, n_777_v);
  spice_node_2 n_n_124(eclk, ereset, n_124_port_5,n_124_port_9, n_124_v);
  spice_node_0 n_n_45(eclk, ereset,  n_45_v);
  spice_node_3 n_db4(eclk, ereset, db4_port_0,db4_port_1,db4_port_3, db4_v);
  spice_node_2 n_n_175(eclk, ereset, n_175_port_3,n_175_port_6, n_175_v);
  spice_node_2 n_n_1225(eclk, ereset, n_1225_port_5,n_1225_port_7, n_1225_v);
  spice_node_4 n_n_181(eclk, ereset, n_181_port_4,n_181_port_5,n_181_port_6,n_181_port_7, n_181_v);
  spice_node_2 n_n_176(eclk, ereset, n_176_port_5,n_176_port_10, n_176_v);
  spice_node_2 n_n_1232(eclk, ereset, n_1232_port_3,n_1232_port_5, n_1232_v);
  spice_node_2 n_n_190(eclk, ereset, n_190_port_0,n_190_port_3, n_190_v);
  spice_node_2 n_n_1218(eclk, ereset, n_1218_port_3,n_1218_port_6, n_1218_v);
  spice_node_2 n_n_1228(eclk, ereset, n_1228_port_5,n_1228_port_7, n_1228_v);
  spice_node_2 n_n_1220(eclk, ereset, n_1220_port_6,n_1220_port_10, n_1220_v);
  spice_node_2 n_n_172(eclk, ereset, n_172_port_4,n_172_port_8, n_172_v);
  spice_node_2 n_n_1168(eclk, ereset, n_1168_port_4,n_1168_port_8, n_1168_v);
  spice_node_2 n_n_1466(eclk, ereset, n_1466_port_3,n_1466_port_4, n_1466_v);
  spice_node_2 n_n_1161(eclk, ereset, n_1161_port_4,n_1161_port_9, n_1161_v);
  spice_node_2 n_n_1051(eclk, ereset, n_1051_port_3,n_1051_port_6, n_1051_v);
  spice_node_2 n_n_75(eclk, ereset, n_75_port_5,n_75_port_6, n_75_v);
  spice_node_2 n_n_77(eclk, ereset, n_77_port_5,n_77_port_8, n_77_v);
  spice_node_2 n_n_1060(eclk, ereset, n_1060_port_3,n_1060_port_5, n_1060_v);
  spice_node_2 n_n_185(eclk, ereset, n_185_port_5,n_185_port_7, n_185_v);
  spice_node_2 n_n_61(eclk, ereset, n_61_port_3,n_61_port_5, n_61_v);
  spice_node_2 n_n_1053(eclk, ereset, n_1053_port_4,n_1053_port_6, n_1053_v);
  spice_node_2 n_n_136(eclk, ereset, n_136_port_5,n_136_port_10, n_136_v);
  spice_node_2 n_n_1221(eclk, ereset, n_1221_port_5,n_1221_port_7, n_1221_v);
  spice_node_1 n__nmi(eclk, ereset, _nmi_port_1, _nmi_v);
  spice_node_2 n_n_56(eclk, ereset, n_56_port_5,n_56_port_11, n_56_v);
  spice_node_2 n_n_1271(eclk, ereset, n_1271_port_4,n_1271_port_6, n_1271_v);
  spice_node_2 n_n_223(eclk, ereset, n_223_port_3,n_223_port_6, n_223_v);
  spice_node_2 n_n_68(eclk, ereset, n_68_port_4,n_68_port_9, n_68_v);
  spice_node_2 n_n_58(eclk, ereset, n_58_port_4,n_58_port_8, n_58_v);
  spice_node_2 n_n_197(eclk, ereset, n_197_port_3,n_197_port_6, n_197_v);
  spice_node_2 n_n_148(eclk, ereset, n_148_port_6,n_148_port_13, n_148_v);
  spice_node_2 n_n_57(eclk, ereset, n_57_port_3,n_57_port_6, n_57_v);
  spice_node_2 n_n_67(eclk, ereset, n_67_port_3,n_67_port_5, n_67_v);
  spice_node_2 n_n_92(eclk, ereset, n_92_port_4,n_92_port_7, n_92_v);
  spice_node_2 n_n_1092(eclk, ereset, n_1092_port_3,n_1092_port_5, n_1092_v);
  spice_node_2 n_n_1043(eclk, ereset, n_1043_port_1,n_1043_port_3, n_1043_v);
  spice_node_2 n_n_1080(eclk, ereset, n_1080_port_4,n_1080_port_8, n_1080_v);
  spice_node_3 n_n_1590(eclk, ereset, n_1590_port_1,n_1590_port_2,n_1590_port_3, n_1590_v);
  spice_node_2 n_n_1095(eclk, ereset, n_1095_port_4,n_1095_port_8, n_1095_v);
  spice_node_2 n_n_120(eclk, ereset, n_120_port_5,n_120_port_9, n_120_v);
  spice_node_2 n_n_1079(eclk, ereset, n_1079_port_3,n_1079_port_5, n_1079_v);
  spice_node_2 n_n_128(eclk, ereset, n_128_port_6,n_128_port_10, n_128_v);
  spice_node_2 n_n_1300(eclk, ereset, n_1300_port_2,n_1300_port_3, n_1300_v);
  spice_node_2 n_n_1302(eclk, ereset, n_1302_port_0,n_1302_port_2, n_1302_v);
  spice_node_2 n_n_1586(eclk, ereset, n_1586_port_4,n_1586_port_6, n_1586_v);
  spice_node_2 n_n_139(eclk, ereset, n_139_port_5,n_139_port_12, n_139_v);
  spice_node_2 n_n_1126(eclk, ereset, n_1126_port_5,n_1126_port_8, n_1126_v);
  spice_node_2 n_n_70(eclk, ereset, n_70_port_4,n_70_port_7, n_70_v);
  spice_node_1 n__busrq(eclk, ereset, _busrq_port_1, _busrq_v);
  spice_node_1 n__wait(eclk, ereset, _wait_port_1, _wait_v);
  spice_node_2 n_n_241(eclk, ereset, n_241_port_5,n_241_port_7, n_241_v);
  spice_node_2 n_n_216(eclk, ereset, n_216_port_5,n_216_port_8, n_216_v);
  spice_node_2 n_n_1320(eclk, ereset, n_1320_port_3,n_1320_port_5, n_1320_v);
  spice_node_2 n_n_240(eclk, ereset, n_240_port_5,n_240_port_8, n_240_v);
  spice_node_2 n_n_214(eclk, ereset, n_214_port_3,n_214_port_5, n_214_v);
  spice_node_2 n_n_150(eclk, ereset, n_150_port_5,n_150_port_11, n_150_v);
  spice_node_2 n_n_1313(eclk, ereset, n_1313_port_3,n_1313_port_6, n_1313_v);
  spice_node_2 n_n_1701(eclk, ereset, n_1701_port_4,n_1701_port_8, n_1701_v);
  spice_node_2 n_ex_dehl0(eclk, ereset, ex_dehl0_port_5,ex_dehl0_port_9, ex_dehl0_v);
  spice_node_2 n_n_1702(eclk, ereset, n_1702_port_4,n_1702_port_8, n_1702_v);
  spice_node_2 n_ex_dehl1(eclk, ereset, ex_dehl1_port_5,ex_dehl1_port_9, ex_dehl1_v);
  spice_node_0 n_n_1709(eclk, ereset,  n_1709_v);
  spice_node_2 n_n_244(eclk, ereset, n_244_port_4,n_244_port_8, n_244_v);
  spice_node_1 n__int(eclk, ereset, _int_port_1, _int_v);
  spice_node_2 n_n_633(eclk, ereset, n_633_port_5,n_633_port_9, n_633_v);
  spice_node_2 n_n_84(eclk, ereset, n_84_port_6,n_84_port_10, n_84_v);
  spice_node_2 n_n_1129(eclk, ereset, n_1129_port_3,n_1129_port_6, n_1129_v);
  spice_node_2 n_ex_af(eclk, ereset, ex_af_port_5,ex_af_port_10, ex_af_v);
  spice_node_4 n_n_647(eclk, ereset, n_647_port_0,n_647_port_3,n_647_port_4,n_647_port_5, n_647_v);
  spice_node_2 n_n_687(eclk, ereset, n_687_port_5,n_687_port_6, n_687_v);
  spice_node_2 n_n_1783(eclk, ereset, n_1783_port_4,n_1783_port_6, n_1783_v);
  spice_node_2 n_n_1773(eclk, ereset, n_1773_port_5,n_1773_port_9, n_1773_v);
  spice_node_2 n_n_89(eclk, ereset, n_89_port_4,n_89_port_5, n_89_v);
  spice_node_1 n_n_689(eclk, ereset, n_689_port_4, n_689_v);
  spice_node_2 n_n_1171(eclk, ereset, n_1171_port_4,n_1171_port_7, n_1171_v);
  spice_node_2 n_n_127(eclk, ereset, n_127_port_3,n_127_port_6, n_127_v);
  spice_node_2 n_n_259(eclk, ereset, n_259_port_5,n_259_port_8, n_259_v);
  spice_node_2 n_n_1341(eclk, ereset, n_1341_port_3,n_1341_port_5, n_1341_v);
  spice_node_2 n_n_1072(eclk, ereset, n_1072_port_5,n_1072_port_7, n_1072_v);
  spice_node_2 n_n_86(eclk, ereset, n_86_port_6,n_86_port_7, n_86_v);
  spice_node_2 n_n_617(eclk, ereset, n_617_port_3,n_617_port_5, n_617_v);
  spice_node_4 n_n_701(eclk, ereset, n_701_port_0,n_701_port_2,n_701_port_3,n_701_port_4, n_701_v);
  spice_node_4 n_n_696(eclk, ereset, n_696_port_1,n_696_port_2,n_696_port_3,n_696_port_4, n_696_v);
  spice_node_3 n_n_1814(eclk, ereset, n_1814_port_1,n_1814_port_2,n_1814_port_3, n_1814_v);
  spice_node_3 n_reg_pcl0(eclk, ereset, reg_pcl0_port_0,reg_pcl0_port_2,reg_pcl0_port_3, reg_pcl0_v);
  spice_node_3 n_n_1815(eclk, ereset, n_1815_port_1,n_1815_port_2,n_1815_port_3, n_1815_v);
  spice_node_3 n_reg_r0(eclk, ereset, reg_r0_port_0,reg_r0_port_2,reg_r0_port_3, reg_r0_v);
  spice_node_3 n_n_1816(eclk, ereset, n_1816_port_1,n_1816_port_2,n_1816_port_3, n_1816_v);
  spice_node_3 n_reg_z0(eclk, ereset, reg_z0_port_0,reg_z0_port_2,reg_z0_port_3, reg_z0_v);
  spice_node_3 n_n_1817(eclk, ereset, n_1817_port_1,n_1817_port_2,n_1817_port_3, n_1817_v);
  spice_node_3 n_reg_spl0(eclk, ereset, reg_spl0_port_0,reg_spl0_port_2,reg_spl0_port_3, reg_spl0_v);
  spice_node_3 n_n_1818(eclk, ereset, n_1818_port_1,n_1818_port_2,n_1818_port_3, n_1818_v);
  spice_node_3 n_reg_iyl0(eclk, ereset, reg_iyl0_port_0,reg_iyl0_port_2,reg_iyl0_port_3, reg_iyl0_v);
  spice_node_3 n_n_1819(eclk, ereset, n_1819_port_1,n_1819_port_2,n_1819_port_3, n_1819_v);
  spice_node_3 n_reg_ixl0(eclk, ereset, reg_ixl0_port_0,reg_ixl0_port_2,reg_ixl0_port_3, reg_ixl0_v);
  spice_node_3 n_n_1820(eclk, ereset, n_1820_port_1,n_1820_port_2,n_1820_port_3, n_1820_v);
  spice_node_3 n_reg_e0(eclk, ereset, reg_e0_port_0,reg_e0_port_2,reg_e0_port_3, reg_e0_v);
  spice_node_3 n_n_1821(eclk, ereset, n_1821_port_1,n_1821_port_2,n_1821_port_3, n_1821_v);
  spice_node_3 n_reg_ee0(eclk, ereset, reg_ee0_port_0,reg_ee0_port_2,reg_ee0_port_3, reg_ee0_v);
  spice_node_3 n_n_1822(eclk, ereset, n_1822_port_1,n_1822_port_2,n_1822_port_3, n_1822_v);
  spice_node_3 n_reg_l0(eclk, ereset, reg_l0_port_0,reg_l0_port_2,reg_l0_port_3, reg_l0_v);
  spice_node_3 n_n_1823(eclk, ereset, n_1823_port_1,n_1823_port_2,n_1823_port_3, n_1823_v);
  spice_node_3 n_reg_ll0(eclk, ereset, reg_ll0_port_0,reg_ll0_port_2,reg_ll0_port_3, reg_ll0_v);
  spice_node_3 n_n_1824(eclk, ereset, n_1824_port_1,n_1824_port_2,n_1824_port_3, n_1824_v);
  spice_node_3 n_reg_c0(eclk, ereset, reg_c0_port_0,reg_c0_port_2,reg_c0_port_3, reg_c0_v);
  spice_node_3 n_n_1825(eclk, ereset, n_1825_port_1,n_1825_port_2,n_1825_port_3, n_1825_v);
  spice_node_3 n_reg_cc0(eclk, ereset, reg_cc0_port_0,reg_cc0_port_2,reg_cc0_port_3, reg_cc0_v);
  spice_node_3 n_n_1826(eclk, ereset, n_1826_port_1,n_1826_port_2,n_1826_port_3, n_1826_v);
  spice_node_3 n_reg_ff0(eclk, ereset, reg_ff0_port_0,reg_ff0_port_2,reg_ff0_port_3, reg_ff0_v);
  spice_node_3 n_n_1827(eclk, ereset, n_1827_port_1,n_1827_port_2,n_1827_port_3, n_1827_v);
  spice_node_3 n_reg_f0(eclk, ereset, reg_f0_port_0,reg_f0_port_2,reg_f0_port_3, reg_f0_v);
  spice_node_14 n_n_708(eclk, ereset, n_708_port_1,n_708_port_4,n_708_port_5,n_708_port_6,n_708_port_7,n_708_port_8,n_708_port_9,n_708_port_10,n_708_port_11,n_708_port_12,n_708_port_13,n_708_port_14,n_708_port_15,n_708_port_17, n_708_v);
  spice_node_3 n_n_709(eclk, ereset, n_709_port_3,n_709_port_4,n_709_port_5, n_709_v);
  spice_node_2 n_n_149(eclk, ereset, n_149_port_5,n_149_port_8, n_149_v);
  spice_node_3 n_n_721(eclk, ereset, n_721_port_2,n_721_port_3,n_721_port_4, n_721_v);
  spice_node_14 n_n_715(eclk, ereset, n_715_port_1,n_715_port_4,n_715_port_5,n_715_port_6,n_715_port_7,n_715_port_8,n_715_port_9,n_715_port_10,n_715_port_11,n_715_port_12,n_715_port_13,n_715_port_14,n_715_port_15,n_715_port_17, n_715_v);
  spice_node_2 n_n_143(eclk, ereset, n_143_port_6,n_143_port_7, n_143_v);
  spice_node_3 n_reg_pcl1(eclk, ereset, reg_pcl1_port_1,reg_pcl1_port_2,reg_pcl1_port_3, reg_pcl1_v);
  spice_node_3 n_n_1890(eclk, ereset, n_1890_port_0,n_1890_port_2,n_1890_port_3, n_1890_v);
  spice_node_3 n_reg_r1(eclk, ereset, reg_r1_port_1,reg_r1_port_2,reg_r1_port_3, reg_r1_v);
  spice_node_3 n_n_1891(eclk, ereset, n_1891_port_0,n_1891_port_2,n_1891_port_3, n_1891_v);
  spice_node_3 n_reg_z1(eclk, ereset, reg_z1_port_1,reg_z1_port_2,reg_z1_port_3, reg_z1_v);
  spice_node_3 n_n_1892(eclk, ereset, n_1892_port_0,n_1892_port_2,n_1892_port_3, n_1892_v);
  spice_node_3 n_reg_spl1(eclk, ereset, reg_spl1_port_1,reg_spl1_port_2,reg_spl1_port_3, reg_spl1_v);
  spice_node_3 n_n_1893(eclk, ereset, n_1893_port_0,n_1893_port_2,n_1893_port_3, n_1893_v);
  spice_node_3 n_reg_iyl1(eclk, ereset, reg_iyl1_port_1,reg_iyl1_port_2,reg_iyl1_port_3, reg_iyl1_v);
  spice_node_3 n_n_1894(eclk, ereset, n_1894_port_0,n_1894_port_2,n_1894_port_3, n_1894_v);
  spice_node_3 n_reg_ixl1(eclk, ereset, reg_ixl1_port_1,reg_ixl1_port_2,reg_ixl1_port_3, reg_ixl1_v);
  spice_node_3 n_n_1895(eclk, ereset, n_1895_port_0,n_1895_port_2,n_1895_port_3, n_1895_v);
  spice_node_3 n_reg_e1(eclk, ereset, reg_e1_port_1,reg_e1_port_2,reg_e1_port_3, reg_e1_v);
  spice_node_3 n_n_1896(eclk, ereset, n_1896_port_0,n_1896_port_2,n_1896_port_3, n_1896_v);
  spice_node_3 n_reg_ee1(eclk, ereset, reg_ee1_port_1,reg_ee1_port_2,reg_ee1_port_3, reg_ee1_v);
  spice_node_3 n_n_1897(eclk, ereset, n_1897_port_0,n_1897_port_2,n_1897_port_3, n_1897_v);
  spice_node_3 n_reg_l1(eclk, ereset, reg_l1_port_1,reg_l1_port_2,reg_l1_port_3, reg_l1_v);
  spice_node_3 n_n_1898(eclk, ereset, n_1898_port_0,n_1898_port_2,n_1898_port_3, n_1898_v);
  spice_node_3 n_reg_ll1(eclk, ereset, reg_ll1_port_1,reg_ll1_port_2,reg_ll1_port_3, reg_ll1_v);
  spice_node_3 n_n_1899(eclk, ereset, n_1899_port_0,n_1899_port_2,n_1899_port_3, n_1899_v);
  spice_node_3 n_reg_c1(eclk, ereset, reg_c1_port_1,reg_c1_port_2,reg_c1_port_3, reg_c1_v);
  spice_node_3 n_n_1900(eclk, ereset, n_1900_port_0,n_1900_port_2,n_1900_port_3, n_1900_v);
  spice_node_3 n_reg_cc1(eclk, ereset, reg_cc1_port_1,reg_cc1_port_2,reg_cc1_port_3, reg_cc1_v);
  spice_node_3 n_n_1901(eclk, ereset, n_1901_port_0,n_1901_port_2,n_1901_port_3, n_1901_v);
  spice_node_3 n_reg_ff1(eclk, ereset, reg_ff1_port_1,reg_ff1_port_2,reg_ff1_port_3, reg_ff1_v);
  spice_node_3 n_n_1902(eclk, ereset, n_1902_port_0,n_1902_port_2,n_1902_port_3, n_1902_v);
  spice_node_3 n_reg_f1(eclk, ereset, reg_f1_port_1,reg_f1_port_2,reg_f1_port_3, reg_f1_v);
  spice_node_3 n_n_1903(eclk, ereset, n_1903_port_0,n_1903_port_2,n_1903_port_3, n_1903_v);
  spice_node_1 n_n_723(eclk, ereset, n_723_port_4, n_723_v);
  spice_node_3 n_n_728(eclk, ereset, n_728_port_2,n_728_port_3,n_728_port_4, n_728_v);
  spice_node_5 n_n_726(eclk, ereset, n_726_port_1,n_726_port_2,n_726_port_3,n_726_port_4,n_726_port_5, n_726_v);
  spice_node_2 n_n_1184(eclk, ereset, n_1184_port_3,n_1184_port_4, n_1184_v);
  spice_node_3 n_n_1915(eclk, ereset, n_1915_port_1,n_1915_port_2,n_1915_port_3, n_1915_v);
  spice_node_3 n_reg_pcl2(eclk, ereset, reg_pcl2_port_0,reg_pcl2_port_2,reg_pcl2_port_3, reg_pcl2_v);
  spice_node_3 n_n_1916(eclk, ereset, n_1916_port_1,n_1916_port_2,n_1916_port_3, n_1916_v);
  spice_node_3 n_reg_r2(eclk, ereset, reg_r2_port_0,reg_r2_port_2,reg_r2_port_3, reg_r2_v);
  spice_node_3 n_n_1917(eclk, ereset, n_1917_port_1,n_1917_port_2,n_1917_port_3, n_1917_v);
  spice_node_3 n_reg_z2(eclk, ereset, reg_z2_port_0,reg_z2_port_2,reg_z2_port_3, reg_z2_v);
  spice_node_3 n_n_1918(eclk, ereset, n_1918_port_1,n_1918_port_2,n_1918_port_3, n_1918_v);
  spice_node_3 n_reg_spl2(eclk, ereset, reg_spl2_port_0,reg_spl2_port_2,reg_spl2_port_3, reg_spl2_v);
  spice_node_3 n_n_1919(eclk, ereset, n_1919_port_1,n_1919_port_2,n_1919_port_3, n_1919_v);
  spice_node_3 n_reg_iyl2(eclk, ereset, reg_iyl2_port_0,reg_iyl2_port_2,reg_iyl2_port_3, reg_iyl2_v);
  spice_node_3 n_n_1920(eclk, ereset, n_1920_port_1,n_1920_port_2,n_1920_port_3, n_1920_v);
  spice_node_3 n_reg_ixl2(eclk, ereset, reg_ixl2_port_0,reg_ixl2_port_2,reg_ixl2_port_3, reg_ixl2_v);
  spice_node_3 n_n_1921(eclk, ereset, n_1921_port_1,n_1921_port_2,n_1921_port_3, n_1921_v);
  spice_node_3 n_reg_e2(eclk, ereset, reg_e2_port_0,reg_e2_port_2,reg_e2_port_3, reg_e2_v);
  spice_node_3 n_n_1922(eclk, ereset, n_1922_port_1,n_1922_port_2,n_1922_port_3, n_1922_v);
  spice_node_3 n_reg_ee2(eclk, ereset, reg_ee2_port_0,reg_ee2_port_2,reg_ee2_port_3, reg_ee2_v);
  spice_node_3 n_n_1923(eclk, ereset, n_1923_port_1,n_1923_port_2,n_1923_port_3, n_1923_v);
  spice_node_3 n_reg_l2(eclk, ereset, reg_l2_port_0,reg_l2_port_2,reg_l2_port_3, reg_l2_v);
  spice_node_3 n_n_1924(eclk, ereset, n_1924_port_1,n_1924_port_2,n_1924_port_3, n_1924_v);
  spice_node_3 n_reg_ll2(eclk, ereset, reg_ll2_port_0,reg_ll2_port_2,reg_ll2_port_3, reg_ll2_v);
  spice_node_3 n_n_1925(eclk, ereset, n_1925_port_1,n_1925_port_2,n_1925_port_3, n_1925_v);
  spice_node_3 n_reg_c2(eclk, ereset, reg_c2_port_0,reg_c2_port_2,reg_c2_port_3, reg_c2_v);
  spice_node_3 n_n_1926(eclk, ereset, n_1926_port_1,n_1926_port_2,n_1926_port_3, n_1926_v);
  spice_node_3 n_reg_cc2(eclk, ereset, reg_cc2_port_0,reg_cc2_port_2,reg_cc2_port_3, reg_cc2_v);
  spice_node_3 n_n_1927(eclk, ereset, n_1927_port_1,n_1927_port_2,n_1927_port_3, n_1927_v);
  spice_node_3 n_reg_ff2(eclk, ereset, reg_ff2_port_0,reg_ff2_port_2,reg_ff2_port_3, reg_ff2_v);
  spice_node_3 n_n_1928(eclk, ereset, n_1928_port_1,n_1928_port_2,n_1928_port_3, n_1928_v);
  spice_node_3 n_reg_f2(eclk, ereset, reg_f2_port_0,reg_f2_port_2,reg_f2_port_3, reg_f2_v);
  spice_node_14 n_n_745(eclk, ereset, n_745_port_1,n_745_port_4,n_745_port_5,n_745_port_6,n_745_port_7,n_745_port_8,n_745_port_9,n_745_port_10,n_745_port_11,n_745_port_12,n_745_port_13,n_745_port_14,n_745_port_15,n_745_port_17, n_745_v);
  spice_node_3 n_n_746(eclk, ereset, n_746_port_3,n_746_port_4,n_746_port_5, n_746_v);
  spice_node_3 n_n_763(eclk, ereset, n_763_port_2,n_763_port_3,n_763_port_4, n_763_v);
  spice_node_14 n_n_753(eclk, ereset, n_753_port_1,n_753_port_2,n_753_port_3,n_753_port_4,n_753_port_5,n_753_port_6,n_753_port_7,n_753_port_8,n_753_port_9,n_753_port_12,n_753_port_13,n_753_port_14,n_753_port_15,n_753_port_17, n_753_v);
  spice_node_3 n_reg_pcl3(eclk, ereset, reg_pcl3_port_1,reg_pcl3_port_2,reg_pcl3_port_3, reg_pcl3_v);
  spice_node_3 n_n_1996(eclk, ereset, n_1996_port_0,n_1996_port_2,n_1996_port_3, n_1996_v);
  spice_node_3 n_reg_r3(eclk, ereset, reg_r3_port_1,reg_r3_port_2,reg_r3_port_3, reg_r3_v);
  spice_node_3 n_n_1997(eclk, ereset, n_1997_port_0,n_1997_port_2,n_1997_port_3, n_1997_v);
  spice_node_3 n_reg_z3(eclk, ereset, reg_z3_port_1,reg_z3_port_2,reg_z3_port_3, reg_z3_v);
  spice_node_3 n_n_1998(eclk, ereset, n_1998_port_0,n_1998_port_2,n_1998_port_3, n_1998_v);
  spice_node_3 n_reg_spl3(eclk, ereset, reg_spl3_port_1,reg_spl3_port_2,reg_spl3_port_3, reg_spl3_v);
  spice_node_3 n_n_1999(eclk, ereset, n_1999_port_0,n_1999_port_2,n_1999_port_3, n_1999_v);
  spice_node_3 n_reg_iyl3(eclk, ereset, reg_iyl3_port_1,reg_iyl3_port_2,reg_iyl3_port_3, reg_iyl3_v);
  spice_node_3 n_n_2000(eclk, ereset, n_2000_port_0,n_2000_port_2,n_2000_port_3, n_2000_v);
  spice_node_3 n_reg_ixl3(eclk, ereset, reg_ixl3_port_1,reg_ixl3_port_2,reg_ixl3_port_3, reg_ixl3_v);
  spice_node_3 n_n_2001(eclk, ereset, n_2001_port_0,n_2001_port_2,n_2001_port_3, n_2001_v);
  spice_node_3 n_reg_e3(eclk, ereset, reg_e3_port_1,reg_e3_port_2,reg_e3_port_3, reg_e3_v);
  spice_node_3 n_n_2002(eclk, ereset, n_2002_port_0,n_2002_port_2,n_2002_port_3, n_2002_v);
  spice_node_3 n_reg_ee3(eclk, ereset, reg_ee3_port_1,reg_ee3_port_2,reg_ee3_port_3, reg_ee3_v);
  spice_node_3 n_n_2003(eclk, ereset, n_2003_port_0,n_2003_port_2,n_2003_port_3, n_2003_v);
  spice_node_3 n_reg_l3(eclk, ereset, reg_l3_port_1,reg_l3_port_2,reg_l3_port_3, reg_l3_v);
  spice_node_3 n_n_2004(eclk, ereset, n_2004_port_0,n_2004_port_2,n_2004_port_3, n_2004_v);
  spice_node_3 n_reg_ll3(eclk, ereset, reg_ll3_port_1,reg_ll3_port_2,reg_ll3_port_3, reg_ll3_v);
  spice_node_3 n_n_2005(eclk, ereset, n_2005_port_0,n_2005_port_2,n_2005_port_3, n_2005_v);
  spice_node_3 n_reg_c3(eclk, ereset, reg_c3_port_1,reg_c3_port_2,reg_c3_port_3, reg_c3_v);
  spice_node_3 n_n_2006(eclk, ereset, n_2006_port_0,n_2006_port_2,n_2006_port_3, n_2006_v);
  spice_node_3 n_reg_cc3(eclk, ereset, reg_cc3_port_1,reg_cc3_port_2,reg_cc3_port_3, reg_cc3_v);
  spice_node_3 n_n_2007(eclk, ereset, n_2007_port_0,n_2007_port_2,n_2007_port_3, n_2007_v);
  spice_node_3 n_reg_ff3(eclk, ereset, reg_ff3_port_1,reg_ff3_port_2,reg_ff3_port_3, reg_ff3_v);
  spice_node_3 n_n_2008(eclk, ereset, n_2008_port_0,n_2008_port_2,n_2008_port_3, n_2008_v);
  spice_node_3 n_reg_f3(eclk, ereset, reg_f3_port_1,reg_f3_port_2,reg_f3_port_3, reg_f3_v);
  spice_node_3 n_n_2009(eclk, ereset, n_2009_port_0,n_2009_port_2,n_2009_port_3, n_2009_v);
  spice_node_2 n_n_94(eclk, ereset, n_94_port_3,n_94_port_6, n_94_v);
  spice_node_3 n_n_2019(eclk, ereset, n_2019_port_1,n_2019_port_2,n_2019_port_3, n_2019_v);
  spice_node_3 n_reg_pcl4(eclk, ereset, reg_pcl4_port_0,reg_pcl4_port_2,reg_pcl4_port_3, reg_pcl4_v);
  spice_node_3 n_n_2020(eclk, ereset, n_2020_port_1,n_2020_port_2,n_2020_port_3, n_2020_v);
  spice_node_3 n_reg_r4(eclk, ereset, reg_r4_port_0,reg_r4_port_2,reg_r4_port_3, reg_r4_v);
  spice_node_3 n_n_2021(eclk, ereset, n_2021_port_1,n_2021_port_2,n_2021_port_3, n_2021_v);
  spice_node_3 n_reg_z4(eclk, ereset, reg_z4_port_0,reg_z4_port_2,reg_z4_port_3, reg_z4_v);
  spice_node_3 n_n_2022(eclk, ereset, n_2022_port_1,n_2022_port_2,n_2022_port_3, n_2022_v);
  spice_node_3 n_reg_spl4(eclk, ereset, reg_spl4_port_0,reg_spl4_port_2,reg_spl4_port_3, reg_spl4_v);
  spice_node_3 n_n_2023(eclk, ereset, n_2023_port_1,n_2023_port_2,n_2023_port_3, n_2023_v);
  spice_node_3 n_reg_iyl4(eclk, ereset, reg_iyl4_port_0,reg_iyl4_port_2,reg_iyl4_port_3, reg_iyl4_v);
  spice_node_3 n_n_2024(eclk, ereset, n_2024_port_1,n_2024_port_2,n_2024_port_3, n_2024_v);
  spice_node_3 n_reg_ixl4(eclk, ereset, reg_ixl4_port_0,reg_ixl4_port_2,reg_ixl4_port_3, reg_ixl4_v);
  spice_node_3 n_n_2025(eclk, ereset, n_2025_port_1,n_2025_port_2,n_2025_port_3, n_2025_v);
  spice_node_3 n_reg_e4(eclk, ereset, reg_e4_port_0,reg_e4_port_2,reg_e4_port_3, reg_e4_v);
  spice_node_3 n_n_2026(eclk, ereset, n_2026_port_1,n_2026_port_2,n_2026_port_3, n_2026_v);
  spice_node_3 n_reg_ee4(eclk, ereset, reg_ee4_port_0,reg_ee4_port_2,reg_ee4_port_3, reg_ee4_v);
  spice_node_3 n_n_2027(eclk, ereset, n_2027_port_1,n_2027_port_2,n_2027_port_3, n_2027_v);
  spice_node_3 n_reg_l4(eclk, ereset, reg_l4_port_0,reg_l4_port_2,reg_l4_port_3, reg_l4_v);
  spice_node_3 n_n_2028(eclk, ereset, n_2028_port_1,n_2028_port_2,n_2028_port_3, n_2028_v);
  spice_node_3 n_reg_ll4(eclk, ereset, reg_ll4_port_0,reg_ll4_port_2,reg_ll4_port_3, reg_ll4_v);
  spice_node_3 n_n_2029(eclk, ereset, n_2029_port_1,n_2029_port_2,n_2029_port_3, n_2029_v);
  spice_node_3 n_reg_c4(eclk, ereset, reg_c4_port_0,reg_c4_port_2,reg_c4_port_3, reg_c4_v);
  spice_node_3 n_n_2030(eclk, ereset, n_2030_port_1,n_2030_port_2,n_2030_port_3, n_2030_v);
  spice_node_3 n_reg_cc4(eclk, ereset, reg_cc4_port_0,reg_cc4_port_2,reg_cc4_port_3, reg_cc4_v);
  spice_node_3 n_n_2031(eclk, ereset, n_2031_port_1,n_2031_port_2,n_2031_port_3, n_2031_v);
  spice_node_3 n_reg_ff4(eclk, ereset, reg_ff4_port_0,reg_ff4_port_2,reg_ff4_port_3, reg_ff4_v);
  spice_node_3 n_n_2032(eclk, ereset, n_2032_port_1,n_2032_port_2,n_2032_port_3, n_2032_v);
  spice_node_3 n_reg_f4(eclk, ereset, reg_f4_port_0,reg_f4_port_2,reg_f4_port_3, reg_f4_v);
  spice_node_14 n_n_785(eclk, ereset, n_785_port_1,n_785_port_4,n_785_port_5,n_785_port_6,n_785_port_7,n_785_port_8,n_785_port_9,n_785_port_10,n_785_port_11,n_785_port_12,n_785_port_13,n_785_port_14,n_785_port_15,n_785_port_17, n_785_v);
  spice_node_3 n_n_787(eclk, ereset, n_787_port_3,n_787_port_4,n_787_port_5, n_787_v);
  spice_node_3 n_n_802(eclk, ereset, n_802_port_2,n_802_port_3,n_802_port_4, n_802_v);
  spice_node_2 n_n_1170(eclk, ereset, n_1170_port_4,n_1170_port_5, n_1170_v);
  spice_node_14 n_n_799(eclk, ereset, n_799_port_1,n_799_port_4,n_799_port_5,n_799_port_6,n_799_port_7,n_799_port_8,n_799_port_9,n_799_port_10,n_799_port_11,n_799_port_12,n_799_port_13,n_799_port_14,n_799_port_15,n_799_port_17, n_799_v);
  spice_node_3 n_reg_pcl5(eclk, ereset, reg_pcl5_port_1,reg_pcl5_port_2,reg_pcl5_port_3, reg_pcl5_v);
  spice_node_3 n_n_2094(eclk, ereset, n_2094_port_0,n_2094_port_2,n_2094_port_3, n_2094_v);
  spice_node_3 n_reg_r5(eclk, ereset, reg_r5_port_1,reg_r5_port_2,reg_r5_port_3, reg_r5_v);
  spice_node_3 n_n_2095(eclk, ereset, n_2095_port_0,n_2095_port_2,n_2095_port_3, n_2095_v);
  spice_node_3 n_reg_z5(eclk, ereset, reg_z5_port_1,reg_z5_port_2,reg_z5_port_3, reg_z5_v);
  spice_node_3 n_n_2096(eclk, ereset, n_2096_port_0,n_2096_port_2,n_2096_port_3, n_2096_v);
  spice_node_3 n_reg_spl5(eclk, ereset, reg_spl5_port_1,reg_spl5_port_2,reg_spl5_port_3, reg_spl5_v);
  spice_node_3 n_n_2097(eclk, ereset, n_2097_port_0,n_2097_port_2,n_2097_port_3, n_2097_v);
  spice_node_3 n_reg_iyl5(eclk, ereset, reg_iyl5_port_1,reg_iyl5_port_2,reg_iyl5_port_3, reg_iyl5_v);
  spice_node_3 n_n_2098(eclk, ereset, n_2098_port_0,n_2098_port_2,n_2098_port_3, n_2098_v);
  spice_node_3 n_reg_ixl5(eclk, ereset, reg_ixl5_port_1,reg_ixl5_port_2,reg_ixl5_port_3, reg_ixl5_v);
  spice_node_3 n_n_2099(eclk, ereset, n_2099_port_0,n_2099_port_2,n_2099_port_3, n_2099_v);
  spice_node_3 n_reg_e5(eclk, ereset, reg_e5_port_1,reg_e5_port_2,reg_e5_port_3, reg_e5_v);
  spice_node_3 n_n_2100(eclk, ereset, n_2100_port_0,n_2100_port_2,n_2100_port_3, n_2100_v);
  spice_node_3 n_reg_ee5(eclk, ereset, reg_ee5_port_1,reg_ee5_port_2,reg_ee5_port_3, reg_ee5_v);
  spice_node_3 n_n_2101(eclk, ereset, n_2101_port_0,n_2101_port_2,n_2101_port_3, n_2101_v);
  spice_node_3 n_reg_l5(eclk, ereset, reg_l5_port_1,reg_l5_port_2,reg_l5_port_3, reg_l5_v);
  spice_node_3 n_n_2102(eclk, ereset, n_2102_port_0,n_2102_port_2,n_2102_port_3, n_2102_v);
  spice_node_3 n_reg_ll5(eclk, ereset, reg_ll5_port_1,reg_ll5_port_2,reg_ll5_port_3, reg_ll5_v);
  spice_node_3 n_n_2103(eclk, ereset, n_2103_port_0,n_2103_port_2,n_2103_port_3, n_2103_v);
  spice_node_3 n_reg_c5(eclk, ereset, reg_c5_port_1,reg_c5_port_2,reg_c5_port_3, reg_c5_v);
  spice_node_3 n_n_2104(eclk, ereset, n_2104_port_0,n_2104_port_2,n_2104_port_3, n_2104_v);
  spice_node_3 n_reg_cc5(eclk, ereset, reg_cc5_port_1,reg_cc5_port_2,reg_cc5_port_3, reg_cc5_v);
  spice_node_3 n_n_2105(eclk, ereset, n_2105_port_0,n_2105_port_2,n_2105_port_3, n_2105_v);
  spice_node_3 n_reg_ff5(eclk, ereset, reg_ff5_port_1,reg_ff5_port_2,reg_ff5_port_3, reg_ff5_v);
  spice_node_3 n_n_2106(eclk, ereset, n_2106_port_0,n_2106_port_2,n_2106_port_3, n_2106_v);
  spice_node_3 n_reg_f5(eclk, ereset, reg_f5_port_1,reg_f5_port_2,reg_f5_port_3, reg_f5_v);
  spice_node_3 n_n_2107(eclk, ereset, n_2107_port_0,n_2107_port_2,n_2107_port_3, n_2107_v);
  spice_node_1 n_n_2116(eclk, ereset, n_2116_port_3, n_2116_v);
  spice_node_2 n_n_359(eclk, ereset, n_359_port_3,n_359_port_6, n_359_v);
  spice_node_3 n_n_2119(eclk, ereset, n_2119_port_1,n_2119_port_2,n_2119_port_3, n_2119_v);
  spice_node_3 n_reg_pcl6(eclk, ereset, reg_pcl6_port_0,reg_pcl6_port_2,reg_pcl6_port_3, reg_pcl6_v);
  spice_node_3 n_n_2120(eclk, ereset, n_2120_port_1,n_2120_port_2,n_2120_port_3, n_2120_v);
  spice_node_3 n_reg_r6(eclk, ereset, reg_r6_port_0,reg_r6_port_2,reg_r6_port_3, reg_r6_v);
  spice_node_3 n_n_2121(eclk, ereset, n_2121_port_1,n_2121_port_2,n_2121_port_3, n_2121_v);
  spice_node_3 n_reg_z6(eclk, ereset, reg_z6_port_0,reg_z6_port_2,reg_z6_port_3, reg_z6_v);
  spice_node_3 n_n_2122(eclk, ereset, n_2122_port_1,n_2122_port_2,n_2122_port_3, n_2122_v);
  spice_node_3 n_reg_spl6(eclk, ereset, reg_spl6_port_0,reg_spl6_port_2,reg_spl6_port_3, reg_spl6_v);
  spice_node_3 n_n_2123(eclk, ereset, n_2123_port_1,n_2123_port_2,n_2123_port_3, n_2123_v);
  spice_node_3 n_reg_iyl6(eclk, ereset, reg_iyl6_port_0,reg_iyl6_port_2,reg_iyl6_port_3, reg_iyl6_v);
  spice_node_3 n_n_2124(eclk, ereset, n_2124_port_1,n_2124_port_2,n_2124_port_3, n_2124_v);
  spice_node_3 n_reg_ixl6(eclk, ereset, reg_ixl6_port_0,reg_ixl6_port_2,reg_ixl6_port_3, reg_ixl6_v);
  spice_node_3 n_n_2125(eclk, ereset, n_2125_port_1,n_2125_port_2,n_2125_port_3, n_2125_v);
  spice_node_3 n_reg_e6(eclk, ereset, reg_e6_port_0,reg_e6_port_2,reg_e6_port_3, reg_e6_v);
  spice_node_3 n_n_2126(eclk, ereset, n_2126_port_1,n_2126_port_2,n_2126_port_3, n_2126_v);
  spice_node_3 n_reg_ee6(eclk, ereset, reg_ee6_port_0,reg_ee6_port_2,reg_ee6_port_3, reg_ee6_v);
  spice_node_3 n_n_2127(eclk, ereset, n_2127_port_1,n_2127_port_2,n_2127_port_3, n_2127_v);
  spice_node_3 n_reg_l6(eclk, ereset, reg_l6_port_0,reg_l6_port_2,reg_l6_port_3, reg_l6_v);
  spice_node_3 n_n_2128(eclk, ereset, n_2128_port_1,n_2128_port_2,n_2128_port_3, n_2128_v);
  spice_node_3 n_reg_ll6(eclk, ereset, reg_ll6_port_0,reg_ll6_port_2,reg_ll6_port_3, reg_ll6_v);
  spice_node_3 n_n_2129(eclk, ereset, n_2129_port_1,n_2129_port_2,n_2129_port_3, n_2129_v);
  spice_node_3 n_reg_c6(eclk, ereset, reg_c6_port_0,reg_c6_port_2,reg_c6_port_3, reg_c6_v);
  spice_node_3 n_n_2130(eclk, ereset, n_2130_port_1,n_2130_port_2,n_2130_port_3, n_2130_v);
  spice_node_3 n_reg_cc6(eclk, ereset, reg_cc6_port_0,reg_cc6_port_2,reg_cc6_port_3, reg_cc6_v);
  spice_node_3 n_n_2131(eclk, ereset, n_2131_port_1,n_2131_port_2,n_2131_port_3, n_2131_v);
  spice_node_3 n_reg_ff6(eclk, ereset, reg_ff6_port_0,reg_ff6_port_2,reg_ff6_port_3, reg_ff6_v);
  spice_node_3 n_n_2132(eclk, ereset, n_2132_port_1,n_2132_port_2,n_2132_port_3, n_2132_v);
  spice_node_3 n_reg_f6(eclk, ereset, reg_f6_port_0,reg_f6_port_2,reg_f6_port_3, reg_f6_v);
  spice_node_14 n_n_834(eclk, ereset, n_834_port_1,n_834_port_4,n_834_port_5,n_834_port_6,n_834_port_7,n_834_port_8,n_834_port_9,n_834_port_10,n_834_port_11,n_834_port_12,n_834_port_13,n_834_port_14,n_834_port_15,n_834_port_17, n_834_v);
  spice_node_3 n_n_835(eclk, ereset, n_835_port_1,n_835_port_2,n_835_port_3, n_835_v);
  spice_node_5 n_n_837(eclk, ereset, n_837_port_1,n_837_port_5,n_837_port_6,n_837_port_8,n_837_port_9, n_837_v);
  spice_node_14 n_n_847(eclk, ereset, n_847_port_1,n_847_port_4,n_847_port_5,n_847_port_6,n_847_port_7,n_847_port_8,n_847_port_9,n_847_port_10,n_847_port_11,n_847_port_12,n_847_port_13,n_847_port_14,n_847_port_15,n_847_port_17, n_847_v);
  spice_node_3 n_n_856(eclk, ereset, n_856_port_3,n_856_port_4,n_856_port_5, n_856_v);
  spice_node_3 n_reg_pcl7(eclk, ereset, reg_pcl7_port_1,reg_pcl7_port_2,reg_pcl7_port_3, reg_pcl7_v);
  spice_node_3 n_n_2196(eclk, ereset, n_2196_port_0,n_2196_port_2,n_2196_port_3, n_2196_v);
  spice_node_3 n_reg_r7(eclk, ereset, reg_r7_port_1,reg_r7_port_2,reg_r7_port_3, reg_r7_v);
  spice_node_3 n_n_2197(eclk, ereset, n_2197_port_0,n_2197_port_2,n_2197_port_3, n_2197_v);
  spice_node_3 n_reg_z7(eclk, ereset, reg_z7_port_1,reg_z7_port_2,reg_z7_port_3, reg_z7_v);
  spice_node_3 n_n_2198(eclk, ereset, n_2198_port_0,n_2198_port_2,n_2198_port_3, n_2198_v);
  spice_node_3 n_reg_spl7(eclk, ereset, reg_spl7_port_1,reg_spl7_port_2,reg_spl7_port_3, reg_spl7_v);
  spice_node_3 n_n_2199(eclk, ereset, n_2199_port_0,n_2199_port_2,n_2199_port_3, n_2199_v);
  spice_node_3 n_reg_iyl7(eclk, ereset, reg_iyl7_port_1,reg_iyl7_port_2,reg_iyl7_port_3, reg_iyl7_v);
  spice_node_3 n_n_2200(eclk, ereset, n_2200_port_0,n_2200_port_2,n_2200_port_3, n_2200_v);
  spice_node_3 n_reg_ixl7(eclk, ereset, reg_ixl7_port_1,reg_ixl7_port_2,reg_ixl7_port_3, reg_ixl7_v);
  spice_node_3 n_n_2201(eclk, ereset, n_2201_port_0,n_2201_port_2,n_2201_port_3, n_2201_v);
  spice_node_3 n_reg_e7(eclk, ereset, reg_e7_port_1,reg_e7_port_2,reg_e7_port_3, reg_e7_v);
  spice_node_3 n_n_2202(eclk, ereset, n_2202_port_0,n_2202_port_2,n_2202_port_3, n_2202_v);
  spice_node_3 n_reg_ee7(eclk, ereset, reg_ee7_port_1,reg_ee7_port_2,reg_ee7_port_3, reg_ee7_v);
  spice_node_3 n_n_2203(eclk, ereset, n_2203_port_0,n_2203_port_2,n_2203_port_3, n_2203_v);
  spice_node_3 n_reg_l7(eclk, ereset, reg_l7_port_1,reg_l7_port_2,reg_l7_port_3, reg_l7_v);
  spice_node_3 n_n_2204(eclk, ereset, n_2204_port_0,n_2204_port_2,n_2204_port_3, n_2204_v);
  spice_node_3 n_reg_ll7(eclk, ereset, reg_ll7_port_1,reg_ll7_port_2,reg_ll7_port_3, reg_ll7_v);
  spice_node_3 n_n_2205(eclk, ereset, n_2205_port_0,n_2205_port_2,n_2205_port_3, n_2205_v);
  spice_node_3 n_reg_c7(eclk, ereset, reg_c7_port_1,reg_c7_port_2,reg_c7_port_3, reg_c7_v);
  spice_node_3 n_n_2206(eclk, ereset, n_2206_port_0,n_2206_port_2,n_2206_port_3, n_2206_v);
  spice_node_3 n_reg_cc7(eclk, ereset, reg_cc7_port_1,reg_cc7_port_2,reg_cc7_port_3, reg_cc7_v);
  spice_node_3 n_n_2207(eclk, ereset, n_2207_port_0,n_2207_port_2,n_2207_port_3, n_2207_v);
  spice_node_3 n_reg_ff7(eclk, ereset, reg_ff7_port_1,reg_ff7_port_2,reg_ff7_port_3, reg_ff7_v);
  spice_node_3 n_n_2208(eclk, ereset, n_2208_port_0,n_2208_port_2,n_2208_port_3, n_2208_v);
  spice_node_3 n_reg_f7(eclk, ereset, reg_f7_port_1,reg_f7_port_2,reg_f7_port_3, reg_f7_v);
  spice_node_3 n_n_2209(eclk, ereset, n_2209_port_0,n_2209_port_2,n_2209_port_3, n_2209_v);
  spice_node_3 n_n_754(eclk, ereset, n_754_port_1,n_754_port_2,n_754_port_5, n_754_v);
  spice_node_4 n_n_867(eclk, ereset, n_867_port_1,n_867_port_3,n_867_port_4,n_867_port_5, n_867_v);
  spice_node_3 n_n_861(eclk, ereset, n_861_port_1,n_861_port_2,n_861_port_3, n_861_v);
  spice_node_3 n_n_2232(eclk, ereset, n_2232_port_1,n_2232_port_2,n_2232_port_3, n_2232_v);
  spice_node_3 n_reg_pch0(eclk, ereset, reg_pch0_port_0,reg_pch0_port_2,reg_pch0_port_3, reg_pch0_v);
  spice_node_3 n_n_2233(eclk, ereset, n_2233_port_1,n_2233_port_2,n_2233_port_3, n_2233_v);
  spice_node_3 n_reg_i0(eclk, ereset, reg_i0_port_0,reg_i0_port_2,reg_i0_port_3, reg_i0_v);
  spice_node_3 n_n_2234(eclk, ereset, n_2234_port_1,n_2234_port_2,n_2234_port_3, n_2234_v);
  spice_node_3 n_reg_w0(eclk, ereset, reg_w0_port_0,reg_w0_port_2,reg_w0_port_3, reg_w0_v);
  spice_node_3 n_n_2235(eclk, ereset, n_2235_port_1,n_2235_port_2,n_2235_port_3, n_2235_v);
  spice_node_3 n_reg_sph0(eclk, ereset, reg_sph0_port_0,reg_sph0_port_2,reg_sph0_port_3, reg_sph0_v);
  spice_node_3 n_n_2236(eclk, ereset, n_2236_port_1,n_2236_port_2,n_2236_port_3, n_2236_v);
  spice_node_3 n_reg_iyh0(eclk, ereset, reg_iyh0_port_0,reg_iyh0_port_2,reg_iyh0_port_3, reg_iyh0_v);
  spice_node_3 n_n_2237(eclk, ereset, n_2237_port_1,n_2237_port_2,n_2237_port_3, n_2237_v);
  spice_node_3 n_reg_ixh0(eclk, ereset, reg_ixh0_port_0,reg_ixh0_port_2,reg_ixh0_port_3, reg_ixh0_v);
  spice_node_3 n_n_2238(eclk, ereset, n_2238_port_1,n_2238_port_2,n_2238_port_3, n_2238_v);
  spice_node_3 n_reg_d0(eclk, ereset, reg_d0_port_0,reg_d0_port_2,reg_d0_port_3, reg_d0_v);
  spice_node_3 n_n_2239(eclk, ereset, n_2239_port_1,n_2239_port_2,n_2239_port_3, n_2239_v);
  spice_node_3 n_reg_dd0(eclk, ereset, reg_dd0_port_0,reg_dd0_port_2,reg_dd0_port_3, reg_dd0_v);
  spice_node_3 n_n_2240(eclk, ereset, n_2240_port_1,n_2240_port_2,n_2240_port_3, n_2240_v);
  spice_node_3 n_reg_h0(eclk, ereset, reg_h0_port_0,reg_h0_port_2,reg_h0_port_3, reg_h0_v);
  spice_node_3 n_n_2241(eclk, ereset, n_2241_port_1,n_2241_port_2,n_2241_port_3, n_2241_v);
  spice_node_3 n_reg_hh0(eclk, ereset, reg_hh0_port_0,reg_hh0_port_2,reg_hh0_port_3, reg_hh0_v);
  spice_node_3 n_n_2242(eclk, ereset, n_2242_port_1,n_2242_port_2,n_2242_port_3, n_2242_v);
  spice_node_3 n_reg_b0(eclk, ereset, reg_b0_port_0,reg_b0_port_2,reg_b0_port_3, reg_b0_v);
  spice_node_3 n_n_2243(eclk, ereset, n_2243_port_1,n_2243_port_2,n_2243_port_3, n_2243_v);
  spice_node_3 n_reg_bb0(eclk, ereset, reg_bb0_port_0,reg_bb0_port_2,reg_bb0_port_3, reg_bb0_v);
  spice_node_3 n_n_2244(eclk, ereset, n_2244_port_1,n_2244_port_2,n_2244_port_3, n_2244_v);
  spice_node_3 n_reg_aa0(eclk, ereset, reg_aa0_port_0,reg_aa0_port_2,reg_aa0_port_3, reg_aa0_v);
  spice_node_3 n_n_2245(eclk, ereset, n_2245_port_1,n_2245_port_2,n_2245_port_3, n_2245_v);
  spice_node_3 n_reg_a0(eclk, ereset, reg_a0_port_0,reg_a0_port_2,reg_a0_port_3, reg_a0_v);
  spice_node_5 n_n_852(eclk, ereset, n_852_port_2,n_852_port_3,n_852_port_5,n_852_port_8,n_852_port_10, n_852_v);
  spice_node_14 n_n_880(eclk, ereset, n_880_port_1,n_880_port_4,n_880_port_5,n_880_port_6,n_880_port_7,n_880_port_8,n_880_port_9,n_880_port_10,n_880_port_11,n_880_port_12,n_880_port_13,n_880_port_14,n_880_port_15,n_880_port_17, n_880_v);
  spice_node_3 n_n_881(eclk, ereset, n_881_port_2,n_881_port_3,n_881_port_4, n_881_v);
  spice_node_2 n_n_1178(eclk, ereset, n_1178_port_3,n_1178_port_6, n_1178_v);
  spice_node_2 n_n_140(eclk, ereset, n_140_port_5,n_140_port_7, n_140_v);
  spice_node_3 n_n_892(eclk, ereset, n_892_port_3,n_892_port_4,n_892_port_5, n_892_v);
  spice_node_14 n_n_886(eclk, ereset, n_886_port_1,n_886_port_4,n_886_port_5,n_886_port_6,n_886_port_7,n_886_port_8,n_886_port_9,n_886_port_10,n_886_port_11,n_886_port_12,n_886_port_13,n_886_port_14,n_886_port_15,n_886_port_17, n_886_v);
  spice_node_3 n_reg_pch1(eclk, ereset, reg_pch1_port_1,reg_pch1_port_2,reg_pch1_port_3, reg_pch1_v);
  spice_node_3 n_n_2306(eclk, ereset, n_2306_port_0,n_2306_port_2,n_2306_port_3, n_2306_v);
  spice_node_3 n_reg_i1(eclk, ereset, reg_i1_port_1,reg_i1_port_2,reg_i1_port_3, reg_i1_v);
  spice_node_3 n_n_2307(eclk, ereset, n_2307_port_0,n_2307_port_2,n_2307_port_3, n_2307_v);
  spice_node_3 n_reg_w1(eclk, ereset, reg_w1_port_1,reg_w1_port_2,reg_w1_port_3, reg_w1_v);
  spice_node_3 n_n_2308(eclk, ereset, n_2308_port_0,n_2308_port_2,n_2308_port_3, n_2308_v);
  spice_node_3 n_reg_sph1(eclk, ereset, reg_sph1_port_1,reg_sph1_port_2,reg_sph1_port_3, reg_sph1_v);
  spice_node_3 n_n_2309(eclk, ereset, n_2309_port_0,n_2309_port_2,n_2309_port_3, n_2309_v);
  spice_node_3 n_reg_iyh1(eclk, ereset, reg_iyh1_port_1,reg_iyh1_port_2,reg_iyh1_port_3, reg_iyh1_v);
  spice_node_3 n_n_2310(eclk, ereset, n_2310_port_0,n_2310_port_2,n_2310_port_3, n_2310_v);
  spice_node_3 n_reg_ixh1(eclk, ereset, reg_ixh1_port_1,reg_ixh1_port_2,reg_ixh1_port_3, reg_ixh1_v);
  spice_node_3 n_n_2311(eclk, ereset, n_2311_port_0,n_2311_port_2,n_2311_port_3, n_2311_v);
  spice_node_3 n_reg_d1(eclk, ereset, reg_d1_port_1,reg_d1_port_2,reg_d1_port_3, reg_d1_v);
  spice_node_3 n_n_2312(eclk, ereset, n_2312_port_0,n_2312_port_2,n_2312_port_3, n_2312_v);
  spice_node_3 n_reg_dd1(eclk, ereset, reg_dd1_port_1,reg_dd1_port_2,reg_dd1_port_3, reg_dd1_v);
  spice_node_3 n_n_2313(eclk, ereset, n_2313_port_0,n_2313_port_2,n_2313_port_3, n_2313_v);
  spice_node_3 n_reg_h1(eclk, ereset, reg_h1_port_1,reg_h1_port_2,reg_h1_port_3, reg_h1_v);
  spice_node_3 n_n_2314(eclk, ereset, n_2314_port_0,n_2314_port_2,n_2314_port_3, n_2314_v);
  spice_node_3 n_reg_hh1(eclk, ereset, reg_hh1_port_1,reg_hh1_port_2,reg_hh1_port_3, reg_hh1_v);
  spice_node_3 n_n_2315(eclk, ereset, n_2315_port_0,n_2315_port_2,n_2315_port_3, n_2315_v);
  spice_node_3 n_reg_b1(eclk, ereset, reg_b1_port_1,reg_b1_port_2,reg_b1_port_3, reg_b1_v);
  spice_node_3 n_n_2316(eclk, ereset, n_2316_port_0,n_2316_port_2,n_2316_port_3, n_2316_v);
  spice_node_3 n_reg_bb1(eclk, ereset, reg_bb1_port_1,reg_bb1_port_2,reg_bb1_port_3, reg_bb1_v);
  spice_node_3 n_n_2317(eclk, ereset, n_2317_port_0,n_2317_port_2,n_2317_port_3, n_2317_v);
  spice_node_3 n_reg_aa1(eclk, ereset, reg_aa1_port_1,reg_aa1_port_2,reg_aa1_port_3, reg_aa1_v);
  spice_node_3 n_n_2318(eclk, ereset, n_2318_port_0,n_2318_port_2,n_2318_port_3, n_2318_v);
  spice_node_3 n_reg_a1(eclk, ereset, reg_a1_port_1,reg_a1_port_2,reg_a1_port_3, reg_a1_v);
  spice_node_3 n_n_2319(eclk, ereset, n_2319_port_0,n_2319_port_2,n_2319_port_3, n_2319_v);
  spice_node_5 n_n_889(eclk, ereset, n_889_port_1,n_889_port_2,n_889_port_3,n_889_port_8,n_889_port_9, n_889_v);
  spice_node_1 n_n_2320(eclk, ereset, n_2320_port_4, n_2320_v);
  spice_node_2 n_n_81(eclk, ereset, n_81_port_6,n_81_port_7, n_81_v);
  spice_node_2 n_n_1076(eclk, ereset, n_1076_port_5,n_1076_port_7, n_1076_v);
  spice_node_3 n_n_2344(eclk, ereset, n_2344_port_1,n_2344_port_2,n_2344_port_3, n_2344_v);
  spice_node_3 n_reg_pch2(eclk, ereset, reg_pch2_port_0,reg_pch2_port_2,reg_pch2_port_3, reg_pch2_v);
  spice_node_3 n_n_2345(eclk, ereset, n_2345_port_1,n_2345_port_2,n_2345_port_3, n_2345_v);
  spice_node_3 n_reg_i2(eclk, ereset, reg_i2_port_0,reg_i2_port_2,reg_i2_port_3, reg_i2_v);
  spice_node_3 n_n_2346(eclk, ereset, n_2346_port_1,n_2346_port_2,n_2346_port_3, n_2346_v);
  spice_node_3 n_reg_w2(eclk, ereset, reg_w2_port_0,reg_w2_port_2,reg_w2_port_3, reg_w2_v);
  spice_node_3 n_n_2347(eclk, ereset, n_2347_port_1,n_2347_port_2,n_2347_port_3, n_2347_v);
  spice_node_3 n_reg_sph2(eclk, ereset, reg_sph2_port_0,reg_sph2_port_2,reg_sph2_port_3, reg_sph2_v);
  spice_node_3 n_n_2348(eclk, ereset, n_2348_port_1,n_2348_port_2,n_2348_port_3, n_2348_v);
  spice_node_3 n_reg_iyh2(eclk, ereset, reg_iyh2_port_0,reg_iyh2_port_2,reg_iyh2_port_3, reg_iyh2_v);
  spice_node_3 n_n_2349(eclk, ereset, n_2349_port_1,n_2349_port_2,n_2349_port_3, n_2349_v);
  spice_node_3 n_reg_ixh2(eclk, ereset, reg_ixh2_port_0,reg_ixh2_port_2,reg_ixh2_port_3, reg_ixh2_v);
  spice_node_3 n_n_2350(eclk, ereset, n_2350_port_1,n_2350_port_2,n_2350_port_3, n_2350_v);
  spice_node_3 n_reg_d2(eclk, ereset, reg_d2_port_0,reg_d2_port_2,reg_d2_port_3, reg_d2_v);
  spice_node_3 n_n_2351(eclk, ereset, n_2351_port_1,n_2351_port_2,n_2351_port_3, n_2351_v);
  spice_node_3 n_reg_dd2(eclk, ereset, reg_dd2_port_0,reg_dd2_port_2,reg_dd2_port_3, reg_dd2_v);
  spice_node_3 n_n_2352(eclk, ereset, n_2352_port_1,n_2352_port_2,n_2352_port_3, n_2352_v);
  spice_node_3 n_reg_h2(eclk, ereset, reg_h2_port_0,reg_h2_port_2,reg_h2_port_3, reg_h2_v);
  spice_node_3 n_n_2353(eclk, ereset, n_2353_port_1,n_2353_port_2,n_2353_port_3, n_2353_v);
  spice_node_3 n_reg_hh2(eclk, ereset, reg_hh2_port_0,reg_hh2_port_2,reg_hh2_port_3, reg_hh2_v);
  spice_node_3 n_n_2354(eclk, ereset, n_2354_port_1,n_2354_port_2,n_2354_port_3, n_2354_v);
  spice_node_3 n_reg_b2(eclk, ereset, reg_b2_port_0,reg_b2_port_2,reg_b2_port_3, reg_b2_v);
  spice_node_3 n_n_2355(eclk, ereset, n_2355_port_1,n_2355_port_2,n_2355_port_3, n_2355_v);
  spice_node_3 n_reg_bb2(eclk, ereset, reg_bb2_port_0,reg_bb2_port_2,reg_bb2_port_3, reg_bb2_v);
  spice_node_3 n_n_2356(eclk, ereset, n_2356_port_1,n_2356_port_2,n_2356_port_3, n_2356_v);
  spice_node_3 n_reg_aa2(eclk, ereset, reg_aa2_port_0,reg_aa2_port_2,reg_aa2_port_3, reg_aa2_v);
  spice_node_3 n_n_2357(eclk, ereset, n_2357_port_1,n_2357_port_2,n_2357_port_3, n_2357_v);
  spice_node_3 n_reg_a2(eclk, ereset, reg_a2_port_0,reg_a2_port_2,reg_a2_port_3, reg_a2_v);
  spice_node_2 n_n_85(eclk, ereset, n_85_port_6,n_85_port_8, n_85_v);
  spice_node_14 n_n_914(eclk, ereset, n_914_port_1,n_914_port_4,n_914_port_5,n_914_port_6,n_914_port_7,n_914_port_8,n_914_port_9,n_914_port_10,n_914_port_11,n_914_port_12,n_914_port_13,n_914_port_14,n_914_port_15,n_914_port_17, n_914_v);
  spice_node_4 n_n_918(eclk, ereset, n_918_port_1,n_918_port_3,n_918_port_4,n_918_port_5, n_918_v);
  spice_node_3 n_n_915(eclk, ereset, n_915_port_2,n_915_port_3,n_915_port_4, n_915_v);
  spice_node_3 n_n_928(eclk, ereset, n_928_port_1,n_928_port_2,n_928_port_3, n_928_v);
  spice_node_2 n_n_157(eclk, ereset, n_157_port_4,n_157_port_8, n_157_v);
  spice_node_14 n_n_923(eclk, ereset, n_923_port_1,n_923_port_4,n_923_port_5,n_923_port_6,n_923_port_7,n_923_port_8,n_923_port_9,n_923_port_10,n_923_port_11,n_923_port_12,n_923_port_13,n_923_port_14,n_923_port_15,n_923_port_17, n_923_v);
  spice_node_3 n_reg_pch3(eclk, ereset, reg_pch3_port_1,reg_pch3_port_2,reg_pch3_port_3, reg_pch3_v);
  spice_node_3 n_n_2429(eclk, ereset, n_2429_port_0,n_2429_port_2,n_2429_port_3, n_2429_v);
  spice_node_3 n_reg_i3(eclk, ereset, reg_i3_port_1,reg_i3_port_2,reg_i3_port_3, reg_i3_v);
  spice_node_3 n_n_2430(eclk, ereset, n_2430_port_0,n_2430_port_2,n_2430_port_3, n_2430_v);
  spice_node_3 n_reg_w3(eclk, ereset, reg_w3_port_1,reg_w3_port_2,reg_w3_port_3, reg_w3_v);
  spice_node_3 n_n_2431(eclk, ereset, n_2431_port_0,n_2431_port_2,n_2431_port_3, n_2431_v);
  spice_node_3 n_reg_sph3(eclk, ereset, reg_sph3_port_1,reg_sph3_port_2,reg_sph3_port_3, reg_sph3_v);
  spice_node_3 n_n_2432(eclk, ereset, n_2432_port_0,n_2432_port_2,n_2432_port_3, n_2432_v);
  spice_node_3 n_reg_iyh3(eclk, ereset, reg_iyh3_port_1,reg_iyh3_port_2,reg_iyh3_port_3, reg_iyh3_v);
  spice_node_3 n_n_2433(eclk, ereset, n_2433_port_0,n_2433_port_2,n_2433_port_3, n_2433_v);
  spice_node_3 n_reg_ixh3(eclk, ereset, reg_ixh3_port_1,reg_ixh3_port_2,reg_ixh3_port_3, reg_ixh3_v);
  spice_node_3 n_n_2434(eclk, ereset, n_2434_port_0,n_2434_port_2,n_2434_port_3, n_2434_v);
  spice_node_3 n_reg_d3(eclk, ereset, reg_d3_port_1,reg_d3_port_2,reg_d3_port_3, reg_d3_v);
  spice_node_3 n_n_2435(eclk, ereset, n_2435_port_0,n_2435_port_2,n_2435_port_3, n_2435_v);
  spice_node_3 n_reg_dd3(eclk, ereset, reg_dd3_port_1,reg_dd3_port_2,reg_dd3_port_3, reg_dd3_v);
  spice_node_3 n_n_2436(eclk, ereset, n_2436_port_0,n_2436_port_2,n_2436_port_3, n_2436_v);
  spice_node_3 n_reg_h3(eclk, ereset, reg_h3_port_1,reg_h3_port_2,reg_h3_port_3, reg_h3_v);
  spice_node_3 n_n_2437(eclk, ereset, n_2437_port_0,n_2437_port_2,n_2437_port_3, n_2437_v);
  spice_node_3 n_reg_hh3(eclk, ereset, reg_hh3_port_1,reg_hh3_port_2,reg_hh3_port_3, reg_hh3_v);
  spice_node_3 n_n_2438(eclk, ereset, n_2438_port_0,n_2438_port_2,n_2438_port_3, n_2438_v);
  spice_node_3 n_reg_b3(eclk, ereset, reg_b3_port_1,reg_b3_port_2,reg_b3_port_3, reg_b3_v);
  spice_node_3 n_n_2439(eclk, ereset, n_2439_port_0,n_2439_port_2,n_2439_port_3, n_2439_v);
  spice_node_3 n_reg_bb3(eclk, ereset, reg_bb3_port_1,reg_bb3_port_2,reg_bb3_port_3, reg_bb3_v);
  spice_node_3 n_n_2440(eclk, ereset, n_2440_port_0,n_2440_port_2,n_2440_port_3, n_2440_v);
  spice_node_3 n_reg_aa3(eclk, ereset, reg_aa3_port_1,reg_aa3_port_2,reg_aa3_port_3, reg_aa3_v);
  spice_node_3 n_n_2441(eclk, ereset, n_2441_port_0,n_2441_port_2,n_2441_port_3, n_2441_v);
  spice_node_3 n_reg_a3(eclk, ereset, reg_a3_port_1,reg_a3_port_2,reg_a3_port_3, reg_a3_v);
  spice_node_3 n_n_2442(eclk, ereset, n_2442_port_0,n_2442_port_2,n_2442_port_3, n_2442_v);
  spice_node_5 n_n_903(eclk, ereset, n_903_port_2,n_903_port_3,n_903_port_5,n_903_port_8,n_903_port_10, n_903_v);
  spice_node_2 n_n_1077(eclk, ereset, n_1077_port_5,n_1077_port_8, n_1077_v);
  spice_node_2 n_n_62(eclk, ereset, n_62_port_3,n_62_port_6, n_62_v);
  spice_node_2 n_n_132(eclk, ereset, n_132_port_3,n_132_port_5, n_132_v);
  spice_node_2 n_n_147(eclk, ereset, n_147_port_4,n_147_port_5, n_147_v);
  spice_node_2 n_n_384(eclk, ereset, n_384_port_3,n_384_port_4, n_384_v);
  spice_node_3 n_n_2450(eclk, ereset, n_2450_port_1,n_2450_port_2,n_2450_port_3, n_2450_v);
  spice_node_3 n_reg_pch4(eclk, ereset, reg_pch4_port_0,reg_pch4_port_2,reg_pch4_port_3, reg_pch4_v);
  spice_node_3 n_n_2451(eclk, ereset, n_2451_port_1,n_2451_port_2,n_2451_port_3, n_2451_v);
  spice_node_3 n_reg_i4(eclk, ereset, reg_i4_port_0,reg_i4_port_2,reg_i4_port_3, reg_i4_v);
  spice_node_3 n_n_2452(eclk, ereset, n_2452_port_1,n_2452_port_2,n_2452_port_3, n_2452_v);
  spice_node_3 n_reg_w4(eclk, ereset, reg_w4_port_0,reg_w4_port_2,reg_w4_port_3, reg_w4_v);
  spice_node_3 n_n_2453(eclk, ereset, n_2453_port_1,n_2453_port_2,n_2453_port_3, n_2453_v);
  spice_node_3 n_reg_sph4(eclk, ereset, reg_sph4_port_0,reg_sph4_port_2,reg_sph4_port_3, reg_sph4_v);
  spice_node_3 n_n_2454(eclk, ereset, n_2454_port_1,n_2454_port_2,n_2454_port_3, n_2454_v);
  spice_node_3 n_reg_iyh4(eclk, ereset, reg_iyh4_port_0,reg_iyh4_port_2,reg_iyh4_port_3, reg_iyh4_v);
  spice_node_3 n_n_2455(eclk, ereset, n_2455_port_1,n_2455_port_2,n_2455_port_3, n_2455_v);
  spice_node_3 n_reg_ixh4(eclk, ereset, reg_ixh4_port_0,reg_ixh4_port_2,reg_ixh4_port_3, reg_ixh4_v);
  spice_node_3 n_n_2456(eclk, ereset, n_2456_port_1,n_2456_port_2,n_2456_port_3, n_2456_v);
  spice_node_3 n_reg_d4(eclk, ereset, reg_d4_port_0,reg_d4_port_2,reg_d4_port_3, reg_d4_v);
  spice_node_3 n_n_2457(eclk, ereset, n_2457_port_1,n_2457_port_2,n_2457_port_3, n_2457_v);
  spice_node_3 n_reg_dd4(eclk, ereset, reg_dd4_port_0,reg_dd4_port_2,reg_dd4_port_3, reg_dd4_v);
  spice_node_3 n_n_2458(eclk, ereset, n_2458_port_1,n_2458_port_2,n_2458_port_3, n_2458_v);
  spice_node_3 n_reg_h4(eclk, ereset, reg_h4_port_0,reg_h4_port_2,reg_h4_port_3, reg_h4_v);
  spice_node_3 n_n_2459(eclk, ereset, n_2459_port_1,n_2459_port_2,n_2459_port_3, n_2459_v);
  spice_node_3 n_reg_hh4(eclk, ereset, reg_hh4_port_0,reg_hh4_port_2,reg_hh4_port_3, reg_hh4_v);
  spice_node_3 n_n_2460(eclk, ereset, n_2460_port_1,n_2460_port_2,n_2460_port_3, n_2460_v);
  spice_node_3 n_reg_b4(eclk, ereset, reg_b4_port_0,reg_b4_port_2,reg_b4_port_3, reg_b4_v);
  spice_node_3 n_n_2461(eclk, ereset, n_2461_port_1,n_2461_port_2,n_2461_port_3, n_2461_v);
  spice_node_3 n_reg_bb4(eclk, ereset, reg_bb4_port_0,reg_bb4_port_2,reg_bb4_port_3, reg_bb4_v);
  spice_node_3 n_n_2462(eclk, ereset, n_2462_port_1,n_2462_port_2,n_2462_port_3, n_2462_v);
  spice_node_3 n_reg_aa4(eclk, ereset, reg_aa4_port_0,reg_aa4_port_2,reg_aa4_port_3, reg_aa4_v);
  spice_node_3 n_n_2463(eclk, ereset, n_2463_port_1,n_2463_port_2,n_2463_port_3, n_2463_v);
  spice_node_3 n_reg_a4(eclk, ereset, reg_a4_port_0,reg_a4_port_2,reg_a4_port_3, reg_a4_v);
  spice_node_5 n_n_937(eclk, ereset, n_937_port_4,n_937_port_5,n_937_port_7,n_937_port_8,n_937_port_9, n_937_v);
  spice_node_2 n_n_98(eclk, ereset, n_98_port_4,n_98_port_8, n_98_v);
  spice_node_3 n_n_950(eclk, ereset, n_950_port_3,n_950_port_4,n_950_port_5, n_950_v);
  spice_node_14 n_n_949(eclk, ereset, n_949_port_1,n_949_port_4,n_949_port_5,n_949_port_6,n_949_port_7,n_949_port_8,n_949_port_9,n_949_port_10,n_949_port_11,n_949_port_12,n_949_port_13,n_949_port_14,n_949_port_15,n_949_port_17, n_949_v);
  spice_node_3 n_n_908(eclk, ereset, n_908_port_1,n_908_port_2,n_908_port_3, n_908_v);
  spice_node_3 n_n_963(eclk, ereset, n_963_port_2,n_963_port_3,n_963_port_4, n_963_v);
  spice_node_14 n_n_959(eclk, ereset, n_959_port_1,n_959_port_4,n_959_port_5,n_959_port_6,n_959_port_7,n_959_port_8,n_959_port_9,n_959_port_10,n_959_port_11,n_959_port_12,n_959_port_13,n_959_port_14,n_959_port_15,n_959_port_17, n_959_v);
  spice_node_3 n_reg_pch5(eclk, ereset, reg_pch5_port_1,reg_pch5_port_2,reg_pch5_port_3, reg_pch5_v);
  spice_node_3 n_n_2539(eclk, ereset, n_2539_port_0,n_2539_port_2,n_2539_port_3, n_2539_v);
  spice_node_3 n_reg_i5(eclk, ereset, reg_i5_port_1,reg_i5_port_2,reg_i5_port_3, reg_i5_v);
  spice_node_3 n_n_2540(eclk, ereset, n_2540_port_0,n_2540_port_2,n_2540_port_3, n_2540_v);
  spice_node_3 n_reg_w5(eclk, ereset, reg_w5_port_1,reg_w5_port_2,reg_w5_port_3, reg_w5_v);
  spice_node_3 n_n_2541(eclk, ereset, n_2541_port_0,n_2541_port_2,n_2541_port_3, n_2541_v);
  spice_node_3 n_reg_sph5(eclk, ereset, reg_sph5_port_1,reg_sph5_port_2,reg_sph5_port_3, reg_sph5_v);
  spice_node_3 n_n_2542(eclk, ereset, n_2542_port_0,n_2542_port_2,n_2542_port_3, n_2542_v);
  spice_node_3 n_reg_iyh5(eclk, ereset, reg_iyh5_port_1,reg_iyh5_port_2,reg_iyh5_port_3, reg_iyh5_v);
  spice_node_3 n_n_2543(eclk, ereset, n_2543_port_0,n_2543_port_2,n_2543_port_3, n_2543_v);
  spice_node_3 n_reg_ixh5(eclk, ereset, reg_ixh5_port_1,reg_ixh5_port_2,reg_ixh5_port_3, reg_ixh5_v);
  spice_node_3 n_n_2544(eclk, ereset, n_2544_port_0,n_2544_port_2,n_2544_port_3, n_2544_v);
  spice_node_3 n_reg_d5(eclk, ereset, reg_d5_port_1,reg_d5_port_2,reg_d5_port_3, reg_d5_v);
  spice_node_3 n_n_2545(eclk, ereset, n_2545_port_0,n_2545_port_2,n_2545_port_3, n_2545_v);
  spice_node_3 n_reg_dd5(eclk, ereset, reg_dd5_port_1,reg_dd5_port_2,reg_dd5_port_3, reg_dd5_v);
  spice_node_3 n_n_2546(eclk, ereset, n_2546_port_0,n_2546_port_2,n_2546_port_3, n_2546_v);
  spice_node_3 n_reg_h5(eclk, ereset, reg_h5_port_1,reg_h5_port_2,reg_h5_port_3, reg_h5_v);
  spice_node_3 n_n_2547(eclk, ereset, n_2547_port_0,n_2547_port_2,n_2547_port_3, n_2547_v);
  spice_node_3 n_reg_hh5(eclk, ereset, reg_hh5_port_1,reg_hh5_port_2,reg_hh5_port_3, reg_hh5_v);
  spice_node_3 n_n_2548(eclk, ereset, n_2548_port_0,n_2548_port_2,n_2548_port_3, n_2548_v);
  spice_node_3 n_reg_b5(eclk, ereset, reg_b5_port_1,reg_b5_port_2,reg_b5_port_3, reg_b5_v);
  spice_node_3 n_n_2549(eclk, ereset, n_2549_port_0,n_2549_port_2,n_2549_port_3, n_2549_v);
  spice_node_3 n_reg_bb5(eclk, ereset, reg_bb5_port_1,reg_bb5_port_2,reg_bb5_port_3, reg_bb5_v);
  spice_node_3 n_n_2550(eclk, ereset, n_2550_port_0,n_2550_port_2,n_2550_port_3, n_2550_v);
  spice_node_3 n_reg_aa5(eclk, ereset, reg_aa5_port_1,reg_aa5_port_2,reg_aa5_port_3, reg_aa5_v);
  spice_node_3 n_n_2551(eclk, ereset, n_2551_port_0,n_2551_port_2,n_2551_port_3, n_2551_v);
  spice_node_3 n_reg_a5(eclk, ereset, reg_a5_port_1,reg_a5_port_2,reg_a5_port_3, reg_a5_v);
  spice_node_3 n_n_2552(eclk, ereset, n_2552_port_0,n_2552_port_2,n_2552_port_3, n_2552_v);
  spice_node_3 n_n_956(eclk, ereset, n_956_port_2,n_956_port_3,n_956_port_4, n_956_v);
  spice_node_5 n_n_951(eclk, ereset, n_951_port_2,n_951_port_3,n_951_port_5,n_951_port_8,n_951_port_10, n_951_v);
  spice_node_3 n_n_2573(eclk, ereset, n_2573_port_1,n_2573_port_2,n_2573_port_3, n_2573_v);
  spice_node_3 n_reg_pch6(eclk, ereset, reg_pch6_port_0,reg_pch6_port_2,reg_pch6_port_3, reg_pch6_v);
  spice_node_3 n_n_2574(eclk, ereset, n_2574_port_1,n_2574_port_2,n_2574_port_3, n_2574_v);
  spice_node_3 n_reg_i6(eclk, ereset, reg_i6_port_0,reg_i6_port_2,reg_i6_port_3, reg_i6_v);
  spice_node_3 n_n_2575(eclk, ereset, n_2575_port_1,n_2575_port_2,n_2575_port_3, n_2575_v);
  spice_node_3 n_reg_w6(eclk, ereset, reg_w6_port_0,reg_w6_port_2,reg_w6_port_3, reg_w6_v);
  spice_node_3 n_n_2576(eclk, ereset, n_2576_port_1,n_2576_port_2,n_2576_port_3, n_2576_v);
  spice_node_3 n_reg_sph6(eclk, ereset, reg_sph6_port_0,reg_sph6_port_2,reg_sph6_port_3, reg_sph6_v);
  spice_node_3 n_n_2577(eclk, ereset, n_2577_port_1,n_2577_port_2,n_2577_port_3, n_2577_v);
  spice_node_3 n_reg_iyh6(eclk, ereset, reg_iyh6_port_0,reg_iyh6_port_2,reg_iyh6_port_3, reg_iyh6_v);
  spice_node_3 n_n_2578(eclk, ereset, n_2578_port_1,n_2578_port_2,n_2578_port_3, n_2578_v);
  spice_node_3 n_reg_ixh6(eclk, ereset, reg_ixh6_port_0,reg_ixh6_port_2,reg_ixh6_port_3, reg_ixh6_v);
  spice_node_3 n_n_2579(eclk, ereset, n_2579_port_1,n_2579_port_2,n_2579_port_3, n_2579_v);
  spice_node_3 n_reg_d6(eclk, ereset, reg_d6_port_0,reg_d6_port_2,reg_d6_port_3, reg_d6_v);
  spice_node_3 n_n_2580(eclk, ereset, n_2580_port_1,n_2580_port_2,n_2580_port_3, n_2580_v);
  spice_node_3 n_reg_dd6(eclk, ereset, reg_dd6_port_0,reg_dd6_port_2,reg_dd6_port_3, reg_dd6_v);
  spice_node_3 n_n_2581(eclk, ereset, n_2581_port_1,n_2581_port_2,n_2581_port_3, n_2581_v);
  spice_node_3 n_reg_h6(eclk, ereset, reg_h6_port_0,reg_h6_port_2,reg_h6_port_3, reg_h6_v);
  spice_node_3 n_n_2582(eclk, ereset, n_2582_port_1,n_2582_port_2,n_2582_port_3, n_2582_v);
  spice_node_3 n_reg_hh6(eclk, ereset, reg_hh6_port_0,reg_hh6_port_2,reg_hh6_port_3, reg_hh6_v);
  spice_node_3 n_n_2583(eclk, ereset, n_2583_port_1,n_2583_port_2,n_2583_port_3, n_2583_v);
  spice_node_3 n_reg_b6(eclk, ereset, reg_b6_port_0,reg_b6_port_2,reg_b6_port_3, reg_b6_v);
  spice_node_3 n_n_2584(eclk, ereset, n_2584_port_1,n_2584_port_2,n_2584_port_3, n_2584_v);
  spice_node_3 n_reg_bb6(eclk, ereset, reg_bb6_port_0,reg_bb6_port_2,reg_bb6_port_3, reg_bb6_v);
  spice_node_3 n_n_2585(eclk, ereset, n_2585_port_1,n_2585_port_2,n_2585_port_3, n_2585_v);
  spice_node_3 n_reg_aa6(eclk, ereset, reg_aa6_port_0,reg_aa6_port_2,reg_aa6_port_3, reg_aa6_v);
  spice_node_3 n_n_2586(eclk, ereset, n_2586_port_1,n_2586_port_2,n_2586_port_3, n_2586_v);
  spice_node_3 n_reg_a6(eclk, ereset, reg_a6_port_0,reg_a6_port_2,reg_a6_port_3, reg_a6_v);
  spice_node_1 n__reset(eclk, ereset, _reset_port_1, _reset_v);
  spice_node_14 n_n_980(eclk, ereset, n_980_port_1,n_980_port_4,n_980_port_5,n_980_port_6,n_980_port_7,n_980_port_8,n_980_port_9,n_980_port_10,n_980_port_11,n_980_port_12,n_980_port_13,n_980_port_14,n_980_port_15,n_980_port_17, n_980_v);
  spice_node_3 n_n_981(eclk, ereset, n_981_port_1,n_981_port_2,n_981_port_3, n_981_v);
  spice_node_1 n_n_2617(eclk, ereset, n_2617_port_4, n_2617_v);
  spice_node_14 n_n_985(eclk, ereset, n_985_port_1,n_985_port_4,n_985_port_5,n_985_port_6,n_985_port_7,n_985_port_8,n_985_port_9,n_985_port_10,n_985_port_11,n_985_port_12,n_985_port_13,n_985_port_14,n_985_port_15,n_985_port_17, n_985_v);
  spice_node_5 n_n_983(eclk, ereset, n_983_port_4,n_983_port_5,n_983_port_7,n_983_port_8,n_983_port_9, n_983_v);
  spice_node_3 n_reg_pch7(eclk, ereset, reg_pch7_port_1,reg_pch7_port_2,reg_pch7_port_3, reg_pch7_v);
  spice_node_3 n_n_2643(eclk, ereset, n_2643_port_0,n_2643_port_2,n_2643_port_3, n_2643_v);
  spice_node_3 n_reg_i7(eclk, ereset, reg_i7_port_1,reg_i7_port_2,reg_i7_port_3, reg_i7_v);
  spice_node_3 n_n_2644(eclk, ereset, n_2644_port_0,n_2644_port_2,n_2644_port_3, n_2644_v);
  spice_node_3 n_reg_w7(eclk, ereset, reg_w7_port_1,reg_w7_port_2,reg_w7_port_3, reg_w7_v);
  spice_node_3 n_n_2645(eclk, ereset, n_2645_port_0,n_2645_port_2,n_2645_port_3, n_2645_v);
  spice_node_3 n_reg_sph7(eclk, ereset, reg_sph7_port_1,reg_sph7_port_2,reg_sph7_port_3, reg_sph7_v);
  spice_node_3 n_n_2646(eclk, ereset, n_2646_port_0,n_2646_port_2,n_2646_port_3, n_2646_v);
  spice_node_3 n_reg_iyh7(eclk, ereset, reg_iyh7_port_1,reg_iyh7_port_2,reg_iyh7_port_3, reg_iyh7_v);
  spice_node_3 n_n_2647(eclk, ereset, n_2647_port_0,n_2647_port_2,n_2647_port_3, n_2647_v);
  spice_node_3 n_reg_ixh7(eclk, ereset, reg_ixh7_port_1,reg_ixh7_port_2,reg_ixh7_port_3, reg_ixh7_v);
  spice_node_3 n_n_2648(eclk, ereset, n_2648_port_0,n_2648_port_2,n_2648_port_3, n_2648_v);
  spice_node_3 n_reg_d7(eclk, ereset, reg_d7_port_1,reg_d7_port_2,reg_d7_port_3, reg_d7_v);
  spice_node_3 n_n_2649(eclk, ereset, n_2649_port_0,n_2649_port_2,n_2649_port_3, n_2649_v);
  spice_node_3 n_reg_dd7(eclk, ereset, reg_dd7_port_1,reg_dd7_port_2,reg_dd7_port_3, reg_dd7_v);
  spice_node_3 n_n_2650(eclk, ereset, n_2650_port_0,n_2650_port_2,n_2650_port_3, n_2650_v);
  spice_node_3 n_reg_h7(eclk, ereset, reg_h7_port_1,reg_h7_port_2,reg_h7_port_3, reg_h7_v);
  spice_node_3 n_n_2651(eclk, ereset, n_2651_port_0,n_2651_port_2,n_2651_port_3, n_2651_v);
  spice_node_3 n_reg_hh7(eclk, ereset, reg_hh7_port_1,reg_hh7_port_2,reg_hh7_port_3, reg_hh7_v);
  spice_node_3 n_n_2652(eclk, ereset, n_2652_port_0,n_2652_port_2,n_2652_port_3, n_2652_v);
  spice_node_3 n_reg_b7(eclk, ereset, reg_b7_port_1,reg_b7_port_2,reg_b7_port_3, reg_b7_v);
  spice_node_3 n_n_2653(eclk, ereset, n_2653_port_0,n_2653_port_2,n_2653_port_3, n_2653_v);
  spice_node_3 n_reg_bb7(eclk, ereset, reg_bb7_port_1,reg_bb7_port_2,reg_bb7_port_3, reg_bb7_v);
  spice_node_3 n_n_2654(eclk, ereset, n_2654_port_0,n_2654_port_2,n_2654_port_3, n_2654_v);
  spice_node_3 n_reg_aa7(eclk, ereset, reg_aa7_port_1,reg_aa7_port_2,reg_aa7_port_3, reg_aa7_v);
  spice_node_3 n_n_2655(eclk, ereset, n_2655_port_0,n_2655_port_2,n_2655_port_3, n_2655_v);
  spice_node_3 n_reg_a7(eclk, ereset, reg_a7_port_1,reg_a7_port_2,reg_a7_port_3, reg_a7_v);
  spice_node_3 n_n_2656(eclk, ereset, n_2656_port_0,n_2656_port_2,n_2656_port_3, n_2656_v);
  spice_node_4 n_n_988(eclk, ereset, n_988_port_1,n_988_port_2,n_988_port_4,n_988_port_5, n_988_v);
  spice_node_3 n_n_1001(eclk, ereset, n_1001_port_2,n_1001_port_3,n_1001_port_4, n_1001_v);
  spice_node_5 n_n_995(eclk, ereset, n_995_port_2,n_995_port_3,n_995_port_4,n_995_port_8,n_995_port_10, n_995_v);
  spice_node_1 n_n_1009(eclk, ereset, n_1009_port_4, n_1009_v);
  spice_node_2 n_n_408(eclk, ereset, n_408_port_4,n_408_port_6, n_408_v);
  spice_node_1 n_n_2700(eclk, ereset, n_2700_port_4, n_2700_v);
  spice_node_1 n_n_2701(eclk, ereset, n_2701_port_4, n_2701_v);
  spice_node_1 n_n_2702(eclk, ereset, n_2702_port_4, n_2702_v);
  spice_node_1 n_n_2703(eclk, ereset, n_2703_port_4, n_2703_v);
  spice_node_1 n_n_2704(eclk, ereset, n_2704_port_4, n_2704_v);
  spice_node_1 n_n_2705(eclk, ereset, n_2705_port_4, n_2705_v);
  spice_node_1 n_n_1014(eclk, ereset, n_1014_port_4, n_1014_v);
  spice_node_1 n_n_1017(eclk, ereset, n_1017_port_4, n_1017_v);
  spice_node_1 n_n_1018(eclk, ereset, n_1018_port_4, n_1018_v);
  spice_node_1 n_n_1020(eclk, ereset, n_1020_port_4, n_1020_v);
  spice_node_2 n_n_118(eclk, ereset, n_118_port_4,n_118_port_7, n_118_v);
  spice_node_2 n_n_169(eclk, ereset, n_169_port_3,n_169_port_6, n_169_v);
  spice_node_2 n_n_1204(eclk, ereset, n_1204_port_3,n_1204_port_5, n_1204_v);
  spice_node_14 n_n_902(eclk, ereset, n_902_port_0,n_902_port_1,n_902_port_2,n_902_port_3,n_902_port_4,n_902_port_5,n_902_port_6,n_902_port_7,n_902_port_8,n_902_port_9,n_902_port_10,n_902_port_11,n_902_port_13,n_902_port_15, n_902_v);
  spice_node_3 n_n_769(eclk, ereset, n_769_port_1,n_769_port_2,n_769_port_3, n_769_v);
  spice_node_14 n_n_906(eclk, ereset, n_906_port_0,n_906_port_1,n_906_port_2,n_906_port_3,n_906_port_4,n_906_port_5,n_906_port_6,n_906_port_7,n_906_port_8,n_906_port_9,n_906_port_10,n_906_port_11,n_906_port_13,n_906_port_15, n_906_v);
  spice_node_2 n_n_1217(eclk, ereset, n_1217_port_2,n_1217_port_4, n_1217_v);
  spice_node_3 n_n_913(eclk, ereset, n_913_port_0,n_913_port_1,n_913_port_3, n_913_v);
  spice_node_2 n_n_328(eclk, ereset, n_328_port_2,n_328_port_3, n_328_v);
  spice_node_14 n_n_775(eclk, ereset, n_775_port_1,n_775_port_3,n_775_port_4,n_775_port_5,n_775_port_6,n_775_port_7,n_775_port_8,n_775_port_9,n_775_port_10,n_775_port_11,n_775_port_12,n_775_port_13,n_775_port_14,n_775_port_15, n_775_v);
  spice_node_0 n_n_1061(eclk, ereset,  n_1061_v);
  spice_node_1 n_n_2775(eclk, ereset, n_2775_port_0, n_2775_v);
  spice_node_1 n_n_2776(eclk, ereset, n_2776_port_0, n_2776_v);
  spice_node_2 n_n_225(eclk, ereset, n_225_port_2,n_225_port_3, n_225_v);
  spice_node_1 n_n_475(eclk, ereset, n_475_port_7, n_475_v);
  spice_node_14 n_n_776(eclk, ereset, n_776_port_0,n_776_port_1,n_776_port_2,n_776_port_3,n_776_port_4,n_776_port_5,n_776_port_6,n_776_port_7,n_776_port_8,n_776_port_9,n_776_port_10,n_776_port_11,n_776_port_13,n_776_port_15, n_776_v);
  spice_node_2 n_n_1383(eclk, ereset, n_1383_port_2,n_1383_port_4, n_1383_v);
  spice_node_3 n_n_784(eclk, ereset, n_784_port_0,n_784_port_1,n_784_port_3, n_784_v);
  spice_node_2 n_n_1090(eclk, ereset, n_1090_port_2,n_1090_port_4, n_1090_v);
  spice_node_3 n_n_929(eclk, ereset, n_929_port_1,n_929_port_2,n_929_port_3, n_929_v);
  spice_node_2 n_n_541(eclk, ereset, n_541_port_2,n_541_port_3, n_541_v);
  spice_node_2 n_n_1405(eclk, ereset, n_1405_port_2,n_1405_port_3, n_1405_v);
  spice_node_2 n_n_1327(eclk, ereset, n_1327_port_2,n_1327_port_3, n_1327_v);
  spice_node_14 n_n_934(eclk, ereset, n_934_port_1,n_934_port_3,n_934_port_4,n_934_port_5,n_934_port_6,n_934_port_7,n_934_port_8,n_934_port_9,n_934_port_10,n_934_port_11,n_934_port_12,n_934_port_13,n_934_port_14,n_934_port_15, n_934_v);
  spice_node_2 n_n_1098(eclk, ereset, n_1098_port_2,n_1098_port_4, n_1098_v);
  spice_node_14 n_n_935(eclk, ereset, n_935_port_0,n_935_port_1,n_935_port_2,n_935_port_3,n_935_port_4,n_935_port_5,n_935_port_6,n_935_port_7,n_935_port_8,n_935_port_9,n_935_port_10,n_935_port_11,n_935_port_13,n_935_port_15, n_935_v);
  spice_node_2 n_n_161(eclk, ereset, n_161_port_2,n_161_port_4, n_161_v);
  spice_node_3 n_n_948(eclk, ereset, n_948_port_0,n_948_port_1,n_948_port_3, n_948_v);
  spice_node_2 n_n_146(eclk, ereset, n_146_port_2,n_146_port_4, n_146_v);
  spice_node_3 n_n_700(eclk, ereset, n_700_port_1,n_700_port_2,n_700_port_3, n_700_v);
  spice_node_3 n_n_804(eclk, ereset, n_804_port_1,n_804_port_2,n_804_port_3, n_804_v);
  spice_node_14 n_n_702(eclk, ereset, n_702_port_0,n_702_port_1,n_702_port_2,n_702_port_3,n_702_port_4,n_702_port_5,n_702_port_6,n_702_port_7,n_702_port_8,n_702_port_9,n_702_port_10,n_702_port_11,n_702_port_13,n_702_port_15, n_702_v);
  spice_node_14 n_n_807(eclk, ereset, n_807_port_1,n_807_port_3,n_807_port_4,n_807_port_5,n_807_port_6,n_807_port_7,n_807_port_8,n_807_port_9,n_807_port_10,n_807_port_11,n_807_port_12,n_807_port_13,n_807_port_14,n_807_port_15, n_807_v);
  spice_node_3 n_n_964(eclk, ereset, n_964_port_1,n_964_port_2,n_964_port_3, n_964_v);
  spice_node_3 n_n_707(eclk, ereset, n_707_port_0,n_707_port_1,n_707_port_3, n_707_v);
  spice_node_14 n_n_809(eclk, ereset, n_809_port_0,n_809_port_1,n_809_port_2,n_809_port_3,n_809_port_4,n_809_port_5,n_809_port_6,n_809_port_7,n_809_port_8,n_809_port_9,n_809_port_10,n_809_port_11,n_809_port_13,n_809_port_15, n_809_v);
  spice_node_3 n_n_833(eclk, ereset, n_833_port_0,n_833_port_1,n_833_port_3, n_833_v);
  spice_node_14 n_n_970(eclk, ereset, n_970_port_1,n_970_port_3,n_970_port_4,n_970_port_5,n_970_port_6,n_970_port_7,n_970_port_8,n_970_port_9,n_970_port_10,n_970_port_11,n_970_port_12,n_970_port_13,n_970_port_14,n_970_port_15, n_970_v);
  spice_node_14 n_n_973(eclk, ereset, n_973_port_0,n_973_port_1,n_973_port_2,n_973_port_3,n_973_port_4,n_973_port_5,n_973_port_6,n_973_port_7,n_973_port_8,n_973_port_9,n_973_port_10,n_973_port_11,n_973_port_13,n_973_port_15, n_973_v);
  spice_node_3 n_n_979(eclk, ereset, n_979_port_0,n_979_port_1,n_979_port_3, n_979_v);
  spice_node_3 n_n_857(eclk, ereset, n_857_port_1,n_857_port_2,n_857_port_3, n_857_v);
  spice_node_2 n_n_1649(eclk, ereset, n_1649_port_2,n_1649_port_4, n_1649_v);
  spice_node_3 n_n_722(eclk, ereset, n_722_port_1,n_722_port_2,n_722_port_3, n_722_v);
  spice_node_3 n_n_994(eclk, ereset, n_994_port_1,n_994_port_2,n_994_port_3, n_994_v);
  spice_node_14 n_n_864(eclk, ereset, n_864_port_1,n_864_port_3,n_864_port_4,n_864_port_5,n_864_port_6,n_864_port_7,n_864_port_8,n_864_port_9,n_864_port_10,n_864_port_11,n_864_port_12,n_864_port_13,n_864_port_14,n_864_port_15, n_864_v);
  spice_node_14 n_n_732(eclk, ereset, n_732_port_1,n_732_port_3,n_732_port_4,n_732_port_5,n_732_port_6,n_732_port_7,n_732_port_8,n_732_port_9,n_732_port_10,n_732_port_11,n_732_port_12,n_732_port_13,n_732_port_14,n_732_port_15, n_732_v);
  spice_node_14 n_n_999(eclk, ereset, n_999_port_1,n_999_port_3,n_999_port_4,n_999_port_5,n_999_port_6,n_999_port_7,n_999_port_8,n_999_port_9,n_999_port_10,n_999_port_11,n_999_port_12,n_999_port_13,n_999_port_14,n_999_port_15, n_999_v);
  spice_node_14 n_n_870(eclk, ereset, n_870_port_0,n_870_port_1,n_870_port_2,n_870_port_3,n_870_port_4,n_870_port_5,n_870_port_6,n_870_port_7,n_870_port_8,n_870_port_9,n_870_port_10,n_870_port_11,n_870_port_13,n_870_port_15, n_870_v);
  spice_node_14 n_n_738(eclk, ereset, n_738_port_0,n_738_port_1,n_738_port_2,n_738_port_3,n_738_port_4,n_738_port_5,n_738_port_6,n_738_port_7,n_738_port_8,n_738_port_9,n_738_port_10,n_738_port_11,n_738_port_13,n_738_port_15, n_738_v);
  spice_node_3 n_n_879(eclk, ereset, n_879_port_0,n_879_port_1,n_879_port_3, n_879_v);
  spice_node_2 n_n_1044(eclk, ereset, n_1044_port_2,n_1044_port_3, n_1044_v);
  spice_node_3 n_n_744(eclk, ereset, n_744_port_0,n_744_port_1,n_744_port_3, n_744_v);
  spice_node_3 n_n_893(eclk, ereset, n_893_port_1,n_893_port_2,n_893_port_3, n_893_v);

endmodule

module spice_node_0(input eclk,ereset, output signed [`W-1:0] v);
  assign v = 0;
endmodule

module spice_node_4(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_2(input eclk,ereset, input signed [`W-1:0] i0,i1, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_3(input eclk,ereset, input signed [`W-1:0] i0,i1,i2, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_6(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_7(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_5(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_1(input eclk,ereset, input signed [`W-1:0] i0, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_14(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11+i12+i13;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_mux_3(input eclk,ereset, input clk0,clk1,clk2, input x0,x1,x2, output reg y);
  wire c0,z0;
  wire c1,z1;
  wire c2,z2;

  assign c0 = clk0;
  assign z0 = x0;

  mux_cascade m0(c0, z0, clk1, x1, c1, z1);
  mux_cascade m1(c1, z1, clk2, x2, c2, z2);

  wire clk = c2;
  wire x = z2;

  always @(posedge eclk)
    if (ereset)
      y <= 0;
    else begin
      if (clk)
        y <= x;
    end

endmodule

module spice_mux_2(input eclk,ereset, input clk0,clk1, input x0,x1, output reg y);
  wire c0,z0;
  wire c1,z1;

  assign c0 = clk0;
  assign z0 = x0;

  mux_cascade m0(c0, z0, clk1, x1, c1, z1);

  wire clk = c1;
  wire x = z1;

  always @(posedge eclk)
    if (ereset)
      y <= 0;
    else begin
      if (clk)
        y <= x;
    end

endmodule

